
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_13_1_1_0_fbd6b6484e0226fdfa7c7e6838ce99f45fe9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:36 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_13_1_1_0
// ------------------------------------------------------------------


module leading_sign_13_1_1_0 (
  mantissa, all_same, rtn
);
  input [12:0] mantissa;
  output all_same;
  output [3:0] rtn;


  // Interconnect Declarations
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire [11:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0;
  wire c_h_1_2;
  wire c_h_1_4;

  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0 = (mantissa[11:0])
      ^ (signext_12_1(~ (mantissa[12])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[9:8]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11:10]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7:6]==2'b11);
  assign c_h_1_2 = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[5:4]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3:2]==2'b11);
  assign c_h_1_4 = c_h_1_2 & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[1:0]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1 &
      c_h_1_4;
  assign all_same = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      = (c_h_1_2 & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3))
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl = ~(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      | (~ c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl = ~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[10:9]!=2'b10))
      & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[6:5]!=2'b10))))
      & c_h_1_2)) & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[2:1]!=2'b10))))
      & c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl
      = ~(MUX_v_2_2_2(({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl}), 2'b11,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4));
  assign rtn = {c_h_1_4 , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl};

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [11:0] signext_12_1;
    input  vector;
  begin
    signext_12_1= {{11{vector}}, vector};
  end
  endfunction

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v5.v 
module mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/leading_sign_18_1_1_0_7b2153b3b691fe1ab68d43c72c494a7b6845_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:37 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_18_1_1_0
// ------------------------------------------------------------------


module leading_sign_18_1_1_0 (
  mantissa, all_same, rtn
);
  input [17:0] mantissa;
  output all_same;
  output [4:0] rtn;


  // Interconnect Declarations
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1;
  wire [16:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_7;

  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0
      = (mantissa[16:0]) ^ (signext_17_1(~ (mantissa[17])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[14:13]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16:15]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12:11]==2'b11);
  assign c_h_1_2 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[10:9]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[6:5]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8:7]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4:3]==2'b11);
  assign c_h_1_5 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[2:1]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[0])
      & c_h_1_7;
  assign all_same = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      = c_h_1_6 & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3))
      & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl
      = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[15:14]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[11:10]!=2'b10))))
      & c_h_1_2)) & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[7:6]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[3:2]!=2'b10))))
      & c_h_1_5)))) & c_h_1_6)) & (~ c_h_1_7)) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign rtn = {c_h_1_7 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl};

  function automatic [16:0] signext_17_1;
    input  vector;
  begin
    signext_17_1= {{16{vector}}, vector};
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Wed Apr 23 22:57:04 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [7:0] fsm_output;
  reg [7:0] fsm_output;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 8'd0,
    main_C_1 = 8'd1,
    main_C_2 = 8'd2,
    main_C_3 = 8'd3,
    main_C_4 = 8'd4,
    main_C_5 = 8'd5,
    main_C_6 = 8'd6,
    main_C_7 = 8'd7,
    main_C_8 = 8'd8,
    main_C_9 = 8'd9,
    main_C_10 = 8'd10,
    main_C_11 = 8'd11,
    main_C_12 = 8'd12,
    main_C_13 = 8'd13,
    main_C_14 = 8'd14,
    main_C_15 = 8'd15,
    main_C_16 = 8'd16,
    main_C_17 = 8'd17,
    main_C_18 = 8'd18,
    main_C_19 = 8'd19,
    main_C_20 = 8'd20,
    main_C_21 = 8'd21,
    main_C_22 = 8'd22,
    main_C_23 = 8'd23,
    main_C_24 = 8'd24,
    main_C_25 = 8'd25,
    main_C_26 = 8'd26,
    main_C_27 = 8'd27,
    main_C_28 = 8'd28,
    main_C_29 = 8'd29,
    main_C_30 = 8'd30,
    main_C_31 = 8'd31,
    main_C_32 = 8'd32,
    main_C_33 = 8'd33,
    main_C_34 = 8'd34,
    main_C_35 = 8'd35,
    main_C_36 = 8'd36,
    main_C_37 = 8'd37,
    main_C_38 = 8'd38,
    main_C_39 = 8'd39,
    main_C_40 = 8'd40,
    main_C_41 = 8'd41,
    main_C_42 = 8'd42,
    main_C_43 = 8'd43,
    main_C_44 = 8'd44,
    main_C_45 = 8'd45,
    main_C_46 = 8'd46,
    main_C_47 = 8'd47,
    main_C_48 = 8'd48,
    main_C_49 = 8'd49,
    main_C_50 = 8'd50,
    main_C_51 = 8'd51,
    main_C_52 = 8'd52,
    main_C_53 = 8'd53,
    main_C_54 = 8'd54,
    main_C_55 = 8'd55,
    main_C_56 = 8'd56,
    main_C_57 = 8'd57,
    main_C_58 = 8'd58,
    main_C_59 = 8'd59,
    main_C_60 = 8'd60,
    main_C_61 = 8'd61,
    main_C_62 = 8'd62,
    main_C_63 = 8'd63,
    main_C_64 = 8'd64,
    main_C_65 = 8'd65,
    main_C_66 = 8'd66,
    main_C_67 = 8'd67,
    main_C_68 = 8'd68,
    main_C_69 = 8'd69,
    main_C_70 = 8'd70,
    main_C_71 = 8'd71,
    main_C_72 = 8'd72,
    main_C_73 = 8'd73,
    main_C_74 = 8'd74,
    main_C_75 = 8'd75,
    main_C_76 = 8'd76,
    main_C_77 = 8'd77,
    main_C_78 = 8'd78,
    main_C_79 = 8'd79,
    main_C_80 = 8'd80,
    main_C_81 = 8'd81,
    main_C_82 = 8'd82,
    main_C_83 = 8'd83,
    main_C_84 = 8'd84,
    main_C_85 = 8'd85,
    main_C_86 = 8'd86,
    main_C_87 = 8'd87,
    main_C_88 = 8'd88,
    main_C_89 = 8'd89,
    main_C_90 = 8'd90,
    main_C_91 = 8'd91,
    main_C_92 = 8'd92,
    main_C_93 = 8'd93,
    main_C_94 = 8'd94,
    main_C_95 = 8'd95,
    main_C_96 = 8'd96,
    main_C_97 = 8'd97,
    main_C_98 = 8'd98,
    main_C_99 = 8'd99,
    main_C_100 = 8'd100,
    main_C_101 = 8'd101,
    main_C_102 = 8'd102,
    main_C_103 = 8'd103,
    main_C_104 = 8'd104,
    main_C_105 = 8'd105,
    main_C_106 = 8'd106,
    main_C_107 = 8'd107,
    main_C_108 = 8'd108,
    main_C_109 = 8'd109,
    main_C_110 = 8'd110,
    main_C_111 = 8'd111,
    main_C_112 = 8'd112,
    main_C_113 = 8'd113,
    main_C_114 = 8'd114,
    main_C_115 = 8'd115,
    main_C_116 = 8'd116,
    main_C_117 = 8'd117,
    main_C_118 = 8'd118,
    main_C_119 = 8'd119,
    main_C_120 = 8'd120,
    main_C_121 = 8'd121,
    main_C_122 = 8'd122,
    main_C_123 = 8'd123,
    main_C_124 = 8'd124,
    main_C_125 = 8'd125,
    main_C_126 = 8'd126,
    main_C_127 = 8'd127,
    main_C_128 = 8'd128,
    main_C_129 = 8'd129,
    main_C_130 = 8'd130;

  reg [7:0] state_var;
  reg [7:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 8'b00000001;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 8'b00000010;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 8'b00000011;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 8'b00000100;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 8'b00000101;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 8'b00000110;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 8'b00000111;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 8'b00001000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 8'b00001001;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 8'b00001010;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 8'b00001011;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 8'b00001100;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 8'b00001101;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 8'b00001110;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 8'b00001111;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 8'b00010000;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 8'b00010001;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 8'b00010010;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 8'b00010011;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 8'b00010100;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 8'b00010101;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 8'b00010110;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 8'b00010111;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 8'b00011000;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 8'b00011001;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 8'b00011010;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 8'b00011011;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 8'b00011100;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 8'b00011101;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 8'b00011110;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 8'b00011111;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 8'b00100000;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 8'b00100001;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 8'b00100010;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 8'b00100011;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 8'b00100100;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 8'b00100101;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 8'b00100110;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 8'b00100111;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 8'b00101000;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 8'b00101001;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 8'b00101010;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 8'b00101011;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 8'b00101100;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 8'b00101101;
        state_var_NS = main_C_46;
      end
      main_C_46 : begin
        fsm_output = 8'b00101110;
        state_var_NS = main_C_47;
      end
      main_C_47 : begin
        fsm_output = 8'b00101111;
        state_var_NS = main_C_48;
      end
      main_C_48 : begin
        fsm_output = 8'b00110000;
        state_var_NS = main_C_49;
      end
      main_C_49 : begin
        fsm_output = 8'b00110001;
        state_var_NS = main_C_50;
      end
      main_C_50 : begin
        fsm_output = 8'b00110010;
        state_var_NS = main_C_51;
      end
      main_C_51 : begin
        fsm_output = 8'b00110011;
        state_var_NS = main_C_52;
      end
      main_C_52 : begin
        fsm_output = 8'b00110100;
        state_var_NS = main_C_53;
      end
      main_C_53 : begin
        fsm_output = 8'b00110101;
        state_var_NS = main_C_54;
      end
      main_C_54 : begin
        fsm_output = 8'b00110110;
        state_var_NS = main_C_55;
      end
      main_C_55 : begin
        fsm_output = 8'b00110111;
        state_var_NS = main_C_56;
      end
      main_C_56 : begin
        fsm_output = 8'b00111000;
        state_var_NS = main_C_57;
      end
      main_C_57 : begin
        fsm_output = 8'b00111001;
        state_var_NS = main_C_58;
      end
      main_C_58 : begin
        fsm_output = 8'b00111010;
        state_var_NS = main_C_59;
      end
      main_C_59 : begin
        fsm_output = 8'b00111011;
        state_var_NS = main_C_60;
      end
      main_C_60 : begin
        fsm_output = 8'b00111100;
        state_var_NS = main_C_61;
      end
      main_C_61 : begin
        fsm_output = 8'b00111101;
        state_var_NS = main_C_62;
      end
      main_C_62 : begin
        fsm_output = 8'b00111110;
        state_var_NS = main_C_63;
      end
      main_C_63 : begin
        fsm_output = 8'b00111111;
        state_var_NS = main_C_64;
      end
      main_C_64 : begin
        fsm_output = 8'b01000000;
        state_var_NS = main_C_65;
      end
      main_C_65 : begin
        fsm_output = 8'b01000001;
        state_var_NS = main_C_66;
      end
      main_C_66 : begin
        fsm_output = 8'b01000010;
        state_var_NS = main_C_67;
      end
      main_C_67 : begin
        fsm_output = 8'b01000011;
        state_var_NS = main_C_68;
      end
      main_C_68 : begin
        fsm_output = 8'b01000100;
        state_var_NS = main_C_69;
      end
      main_C_69 : begin
        fsm_output = 8'b01000101;
        state_var_NS = main_C_70;
      end
      main_C_70 : begin
        fsm_output = 8'b01000110;
        state_var_NS = main_C_71;
      end
      main_C_71 : begin
        fsm_output = 8'b01000111;
        state_var_NS = main_C_72;
      end
      main_C_72 : begin
        fsm_output = 8'b01001000;
        state_var_NS = main_C_73;
      end
      main_C_73 : begin
        fsm_output = 8'b01001001;
        state_var_NS = main_C_74;
      end
      main_C_74 : begin
        fsm_output = 8'b01001010;
        state_var_NS = main_C_75;
      end
      main_C_75 : begin
        fsm_output = 8'b01001011;
        state_var_NS = main_C_76;
      end
      main_C_76 : begin
        fsm_output = 8'b01001100;
        state_var_NS = main_C_77;
      end
      main_C_77 : begin
        fsm_output = 8'b01001101;
        state_var_NS = main_C_78;
      end
      main_C_78 : begin
        fsm_output = 8'b01001110;
        state_var_NS = main_C_79;
      end
      main_C_79 : begin
        fsm_output = 8'b01001111;
        state_var_NS = main_C_80;
      end
      main_C_80 : begin
        fsm_output = 8'b01010000;
        state_var_NS = main_C_81;
      end
      main_C_81 : begin
        fsm_output = 8'b01010001;
        state_var_NS = main_C_82;
      end
      main_C_82 : begin
        fsm_output = 8'b01010010;
        state_var_NS = main_C_83;
      end
      main_C_83 : begin
        fsm_output = 8'b01010011;
        state_var_NS = main_C_84;
      end
      main_C_84 : begin
        fsm_output = 8'b01010100;
        state_var_NS = main_C_85;
      end
      main_C_85 : begin
        fsm_output = 8'b01010101;
        state_var_NS = main_C_86;
      end
      main_C_86 : begin
        fsm_output = 8'b01010110;
        state_var_NS = main_C_87;
      end
      main_C_87 : begin
        fsm_output = 8'b01010111;
        state_var_NS = main_C_88;
      end
      main_C_88 : begin
        fsm_output = 8'b01011000;
        state_var_NS = main_C_89;
      end
      main_C_89 : begin
        fsm_output = 8'b01011001;
        state_var_NS = main_C_90;
      end
      main_C_90 : begin
        fsm_output = 8'b01011010;
        state_var_NS = main_C_91;
      end
      main_C_91 : begin
        fsm_output = 8'b01011011;
        state_var_NS = main_C_92;
      end
      main_C_92 : begin
        fsm_output = 8'b01011100;
        state_var_NS = main_C_93;
      end
      main_C_93 : begin
        fsm_output = 8'b01011101;
        state_var_NS = main_C_94;
      end
      main_C_94 : begin
        fsm_output = 8'b01011110;
        state_var_NS = main_C_95;
      end
      main_C_95 : begin
        fsm_output = 8'b01011111;
        state_var_NS = main_C_96;
      end
      main_C_96 : begin
        fsm_output = 8'b01100000;
        state_var_NS = main_C_97;
      end
      main_C_97 : begin
        fsm_output = 8'b01100001;
        state_var_NS = main_C_98;
      end
      main_C_98 : begin
        fsm_output = 8'b01100010;
        state_var_NS = main_C_99;
      end
      main_C_99 : begin
        fsm_output = 8'b01100011;
        state_var_NS = main_C_100;
      end
      main_C_100 : begin
        fsm_output = 8'b01100100;
        state_var_NS = main_C_101;
      end
      main_C_101 : begin
        fsm_output = 8'b01100101;
        state_var_NS = main_C_102;
      end
      main_C_102 : begin
        fsm_output = 8'b01100110;
        state_var_NS = main_C_103;
      end
      main_C_103 : begin
        fsm_output = 8'b01100111;
        state_var_NS = main_C_104;
      end
      main_C_104 : begin
        fsm_output = 8'b01101000;
        state_var_NS = main_C_105;
      end
      main_C_105 : begin
        fsm_output = 8'b01101001;
        state_var_NS = main_C_106;
      end
      main_C_106 : begin
        fsm_output = 8'b01101010;
        state_var_NS = main_C_107;
      end
      main_C_107 : begin
        fsm_output = 8'b01101011;
        state_var_NS = main_C_108;
      end
      main_C_108 : begin
        fsm_output = 8'b01101100;
        state_var_NS = main_C_109;
      end
      main_C_109 : begin
        fsm_output = 8'b01101101;
        state_var_NS = main_C_110;
      end
      main_C_110 : begin
        fsm_output = 8'b01101110;
        state_var_NS = main_C_111;
      end
      main_C_111 : begin
        fsm_output = 8'b01101111;
        state_var_NS = main_C_112;
      end
      main_C_112 : begin
        fsm_output = 8'b01110000;
        state_var_NS = main_C_113;
      end
      main_C_113 : begin
        fsm_output = 8'b01110001;
        state_var_NS = main_C_114;
      end
      main_C_114 : begin
        fsm_output = 8'b01110010;
        state_var_NS = main_C_115;
      end
      main_C_115 : begin
        fsm_output = 8'b01110011;
        state_var_NS = main_C_116;
      end
      main_C_116 : begin
        fsm_output = 8'b01110100;
        state_var_NS = main_C_117;
      end
      main_C_117 : begin
        fsm_output = 8'b01110101;
        state_var_NS = main_C_118;
      end
      main_C_118 : begin
        fsm_output = 8'b01110110;
        state_var_NS = main_C_119;
      end
      main_C_119 : begin
        fsm_output = 8'b01110111;
        state_var_NS = main_C_120;
      end
      main_C_120 : begin
        fsm_output = 8'b01111000;
        state_var_NS = main_C_121;
      end
      main_C_121 : begin
        fsm_output = 8'b01111001;
        state_var_NS = main_C_122;
      end
      main_C_122 : begin
        fsm_output = 8'b01111010;
        state_var_NS = main_C_123;
      end
      main_C_123 : begin
        fsm_output = 8'b01111011;
        state_var_NS = main_C_124;
      end
      main_C_124 : begin
        fsm_output = 8'b01111100;
        state_var_NS = main_C_125;
      end
      main_C_125 : begin
        fsm_output = 8'b01111101;
        state_var_NS = main_C_126;
      end
      main_C_126 : begin
        fsm_output = 8'b01111110;
        state_var_NS = main_C_127;
      end
      main_C_127 : begin
        fsm_output = 8'b01111111;
        state_var_NS = main_C_128;
      end
      main_C_128 : begin
        fsm_output = 8'b10000000;
        state_var_NS = main_C_129;
      end
      main_C_129 : begin
        fsm_output = 8'b10000001;
        state_var_NS = main_C_130;
      end
      main_C_130 : begin
        fsm_output = 8'b10000010;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 8'b00000000;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core_wait_dp
// ------------------------------------------------------------------


module fir_core_wait_dp (
  clk, rst, MAC_1_leading_sign_18_1_1_0_cmp_all_same, MAC_1_leading_sign_18_1_1_0_cmp_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg
);
  input clk;
  input rst;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  output MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;


  // Interconnect Declarations
  reg MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;


  // Interconnect Declarations for Component Instantiations 
  assign MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= 5'b00000;
    end
    else begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, input_m_rsc_dat, input_m_triosy_lz, input_e_rsc_dat, input_e_triosy_lz,
      taps_m_rsc_dat, taps_m_triosy_lz, taps_e_rsc_dat, taps_e_triosy_lz, return_m_rsc_dat,
      return_m_triosy_lz, return_e_rsc_dat, return_e_triosy_lz, MAC_1_leading_sign_18_1_1_0_cmp_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_all_same, MAC_1_leading_sign_18_1_1_0_cmp_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_1_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn, MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_3_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn, MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_5_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn, MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_7_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn, MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_9_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn, MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_11_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn, MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_13_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn, MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_15_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn, MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_17_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn, MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_19_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn, MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_21_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn, MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_23_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn, MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_25_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn, MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_27_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn, MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_29_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn, MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_31_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn
);
  input clk;
  input rst;
  input [10:0] input_m_rsc_dat;
  output input_m_triosy_lz;
  input [4:0] input_e_rsc_dat;
  output input_e_triosy_lz;
  input [351:0] taps_m_rsc_dat;
  output taps_m_triosy_lz;
  input [159:0] taps_e_rsc_dat;
  output taps_e_triosy_lz;
  output [10:0] return_m_rsc_dat;
  output return_m_triosy_lz;
  output [4:0] return_e_rsc_dat;
  output return_e_triosy_lz;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;


  // Interconnect Declarations
  wire [10:0] input_m_rsci_idat;
  wire [4:0] input_e_rsci_idat;
  wire [351:0] taps_m_rsci_idat;
  wire [159:0] taps_e_rsci_idat;
  reg [10:0] return_m_rsci_idat;
  reg [4:0] return_e_rsci_idat;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  wire [7:0] fsm_output;
  wire [5:0] MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_3_result_operator_result_operator_nor_tmp;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp;
  wire [5:0] MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp;
  wire [2:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp;
  wire [2:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire or_tmp_1;
  wire or_tmp_2;
  wire and_dcpl_1;
  wire or_tmp_17;
  wire nor_tmp_9;
  wire or_tmp_25;
  wire and_tmp_3;
  wire nor_tmp_12;
  wire mux_tmp_73;
  wire or_tmp_62;
  wire or_tmp_87;
  wire and_dcpl_36;
  wire or_dcpl_50;
  wire or_dcpl_54;
  wire or_dcpl_56;
  wire and_dcpl_47;
  wire and_dcpl_48;
  wire and_dcpl_49;
  wire and_dcpl_50;
  wire and_dcpl_59;
  wire and_dcpl_60;
  wire and_dcpl_61;
  wire and_dcpl_63;
  wire and_dcpl_64;
  wire and_dcpl_65;
  wire and_dcpl_66;
  wire and_dcpl_67;
  wire mux_tmp_110;
  wire or_tmp_92;
  wire mux_tmp_113;
  wire mux_tmp_116;
  wire not_tmp_115;
  wire mux_tmp_119;
  wire or_tmp_96;
  wire or_tmp_100;
  wire nor_tmp_24;
  wire mux_tmp_126;
  wire or_dcpl_66;
  wire or_tmp_102;
  wire mux_tmp_128;
  wire mux_tmp_129;
  wire and_tmp_6;
  wire mux_tmp_131;
  wire and_tmp_7;
  wire and_tmp_8;
  wire or_tmp_104;
  wire or_tmp_105;
  wire mux_tmp_136;
  wire mux_tmp_138;
  wire or_dcpl_68;
  wire or_dcpl_71;
  wire and_dcpl_89;
  wire and_dcpl_90;
  wire and_dcpl_91;
  wire and_dcpl_93;
  wire and_dcpl_95;
  wire and_dcpl_96;
  wire or_dcpl_74;
  wire or_dcpl_75;
  wire and_dcpl_98;
  wire and_dcpl_99;
  wire and_dcpl_100;
  wire and_dcpl_101;
  wire xor_dcpl_3;
  wire and_dcpl_103;
  wire and_dcpl_104;
  wire nor_tmp_27;
  wire or_tmp_110;
  wire mux_tmp_145;
  wire not_tmp_131;
  wire mux_tmp_147;
  wire mux_tmp_149;
  wire mux_tmp_151;
  wire and_tmp_9;
  wire and_tmp_10;
  wire and_tmp_11;
  wire or_tmp_114;
  wire and_dcpl_118;
  wire or_tmp_116;
  wire or_dcpl_83;
  wire nor_tmp_29;
  wire and_dcpl_129;
  wire and_dcpl_132;
  wire and_dcpl_135;
  wire and_dcpl_136;
  wire and_dcpl_143;
  wire and_dcpl_148;
  wire or_dcpl_89;
  wire or_dcpl_96;
  wire and_dcpl_167;
  wire or_dcpl_100;
  wire or_tmp_128;
  wire and_dcpl_290;
  wire mux_tmp_201;
  wire and_dcpl_323;
  wire and_dcpl_324;
  wire and_dcpl_341;
  wire and_dcpl_343;
  wire and_dcpl_347;
  wire and_dcpl_354;
  wire and_dcpl_355;
  wire and_dcpl_360;
  wire and_dcpl_365;
  wire and_dcpl_382;
  wire and_dcpl_399;
  wire and_dcpl_416;
  wire and_dcpl_417;
  wire and_dcpl_422;
  wire and_dcpl_427;
  wire and_dcpl_432;
  wire or_tmp_204;
  wire or_dcpl_170;
  wire mux_tmp_284;
  wire mux_tmp_285;
  wire and_dcpl_505;
  wire and_dcpl_514;
  wire and_dcpl_518;
  wire and_dcpl_524;
  wire and_dcpl_529;
  wire and_dcpl_533;
  wire and_dcpl_543;
  wire and_dcpl_547;
  wire and_dcpl_557;
  wire and_dcpl_558;
  wire and_dcpl_564;
  wire and_dcpl_569;
  wire and_dcpl_570;
  wire and_dcpl_574;
  wire and_dcpl_578;
  wire and_dcpl_587;
  wire and_dcpl_589;
  wire and_dcpl_593;
  wire and_dcpl_609;
  wire and_dcpl_613;
  wire not_tmp_342;
  wire or_dcpl_180;
  wire nor_tmp_33;
  wire nor_tmp_36;
  wire mux_tmp_351;
  wire or_dcpl_200;
  wire and_dcpl_688;
  wire and_dcpl_724;
  reg ac_float_cctor_operator_return_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  reg ac_float_cctor_operator_return_9_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  reg result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  wire [10:0] MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1;
  wire MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w1;
  wire MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w1;
  wire MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w1;
  wire MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w1;
  wire MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w1;
  wire MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w1;
  wire MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2;
  wire MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2;
  wire MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2;
  wire MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2;
  wire MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2;
  wire MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2;
  wire MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2;
  wire MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva;
  reg MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva;
  reg MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva;
  reg MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva;
  reg MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva;
  reg MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva;
  reg MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva;
  reg MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva;
  reg MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva;
  reg MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva;
  reg MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva;
  reg MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva;
  reg MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva;
  reg MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva;
  reg MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva;
  reg MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva;
  reg MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  reg [10:0] delay_lane_m_30_sva;
  reg [10:0] delay_lane_m_29_sva;
  reg [10:0] delay_lane_m_28_sva;
  reg [10:0] delay_lane_m_27_sva;
  reg [10:0] delay_lane_m_26_sva;
  reg [10:0] delay_lane_m_25_sva;
  reg [10:0] delay_lane_m_24_sva;
  reg [10:0] delay_lane_m_23_sva;
  reg [10:0] delay_lane_m_22_sva;
  reg [10:0] delay_lane_m_21_sva;
  reg [10:0] delay_lane_m_20_sva;
  reg [10:0] delay_lane_m_19_sva;
  reg [10:0] delay_lane_m_18_sva;
  reg [10:0] delay_lane_m_17_sva;
  reg [10:0] delay_lane_m_16_sva;
  reg [10:0] delay_lane_m_15_sva;
  reg [10:0] delay_lane_m_14_sva;
  reg [10:0] delay_lane_m_13_sva;
  reg [10:0] delay_lane_m_12_sva;
  reg [10:0] delay_lane_m_11_sva;
  reg [10:0] delay_lane_m_10_sva;
  reg [10:0] delay_lane_m_9_sva;
  reg [10:0] delay_lane_m_8_sva;
  reg [10:0] delay_lane_m_7_sva;
  reg [10:0] delay_lane_m_6_sva;
  reg [10:0] delay_lane_m_5_sva;
  reg [10:0] delay_lane_m_4_sva;
  reg [10:0] delay_lane_m_3_sva;
  reg [10:0] delay_lane_m_1_sva;
  reg [10:0] delay_lane_m_0_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
  wire [6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_seb;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0;
  wire [6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_seb;
  wire and_135_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0;
  wire [6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_seb;
  wire and_134_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0;
  wire [6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_seb;
  wire and_133_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0;
  wire [6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_seb;
  wire and_132_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0;
  wire [6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_seb;
  wire and_131_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0;
  wire [6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_seb;
  wire and_129_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0;
  wire [6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_seb;
  wire nor_113_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0;
  wire [6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_seb;
  wire nor_112_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0;
  wire [6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_seb;
  wire nor_111_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0;
  wire [6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_seb;
  wire nor_110_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0;
  wire [6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_seb;
  wire nor_109_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0;
  wire [6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_seb;
  wire nor_108_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0;
  wire [6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_seb;
  wire nor_107_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0;
  wire [6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_seb;
  wire nor_106_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_ssc;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse;
  wire or_138_cse;
  wire nor_179_cse;
  wire or_359_cse;
  wire or_165_cse;
  wire nor_160_cse;
  reg reg_return_e_triosy_obj_ld_cse;
  reg reg_taps_e_triosy_obj_ld_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse;
  wire nor_202_cse;
  wire nor_231_cse;
  wire nor_227_cse;
  wire nor_223_cse;
  wire nor_219_cse;
  wire nor_214_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse;
  wire or_183_cse;
  wire nor_187_cse;
  wire nor_190_cse;
  wire nor_193_cse;
  wire nor_196_cse;
  wire nor_199_cse;
  wire nor_207_cse;
  wire nor_210_cse;
  wire nor_212_cse;
  wire nor_177_cse;
  wire nor_175_cse;
  wire nor_173_cse;
  wire nor_166_cse;
  wire nor_164_cse;
  wire nor_169_cse;
  wire nor_61_cse;
  wire nor_66_cse;
  wire and_867_cse;
  wire and_861_cse;
  wire and_880_cse;
  wire nor_203_cse;
  wire or_495_cse;
  wire or_92_cse;
  wire mux_420_cse;
  wire mux_419_cse;
  wire mux_416_cse;
  wire mux_409_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc;
  reg [3:0] MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0;
  reg [3:0] MAC_ac_float_cctor_m_4_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0;
  reg MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5;
  wire or_tmp_270;
  wire and_tmp_15;
  wire or_tmp_283;
  wire or_tmp_294;
  wire mux_tmp_427;
  wire nor_tmp_73;
  wire mux_tmp_434;
  wire mux_tmp_435;
  wire mux_tmp_436;
  wire mux_tmp_437;
  wire mux_tmp_438;
  wire mux_tmp_439;
  wire mux_tmp_440;
  wire mux_tmp_441;
  wire mux_tmp_442;
  wire mux_tmp_445;
  wire mux_tmp_448;
  wire mux_tmp_451;
  wire mux_tmp_454;
  reg [6:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0;
  wire or_553_tmp;
  wire and_698_m1c;
  wire and_703_m1c;
  wire and_704_m1c;
  wire and_705_m1c;
  wire and_706_m1c;
  wire and_707_m1c;
  wire and_708_m1c;
  wire and_709_m1c;
  wire and_710_m1c;
  wire and_711_m1c;
  wire and_712_m1c;
  wire and_713_m1c;
  wire and_714_m1c;
  wire and_715_m1c;
  wire and_716_m1c;
  wire and_717_m1c;
  wire and_718_m1c;
  wire and_719_m1c;
  wire and_720_m1c;
  wire and_721_m1c;
  wire and_722_m1c;
  wire and_723_m1c;
  wire and_724_m1c;
  wire and_725_m1c;
  wire and_726_m1c;
  wire and_727_m1c;
  wire and_728_m1c;
  wire and_729_m1c;
  wire and_730_m1c;
  wire and_731_m1c;
  wire and_732_m1c;
  wire mux_461_tmp;
  wire and_929_cse;
  wire and_899_cse;
  wire and_902_cse;
  wire [5:0] MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [12:0] MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [11:0] MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [12:0] MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] z_out;
  wire [12:0] z_out_1;
  wire [12:0] z_out_2;
  wire [12:0] z_out_3;
  wire [12:0] z_out_4;
  wire [12:0] z_out_5;
  wire [12:0] z_out_6;
  wire [12:0] z_out_7;
  wire [12:0] z_out_8;
  wire [12:0] z_out_9;
  wire [12:0] z_out_10;
  wire [12:0] z_out_11;
  wire [12:0] z_out_12;
  wire [12:0] z_out_13;
  wire [12:0] z_out_14;
  wire [6:0] z_out_15;
  wire [5:0] z_out_16;
  wire [6:0] nl_z_out_16;
  wire [10:0] z_out_17;
  reg [10:0] delay_lane_m_2_sva;
  reg [4:0] delay_lane_e_15_sva;
  reg [4:0] delay_lane_e_16_sva;
  reg [4:0] delay_lane_e_14_sva;
  reg [4:0] delay_lane_e_17_sva;
  reg [4:0] delay_lane_e_13_sva;
  reg [4:0] delay_lane_e_18_sva;
  reg [4:0] delay_lane_e_12_sva;
  reg [4:0] delay_lane_e_19_sva;
  reg [4:0] delay_lane_e_11_sva;
  reg [4:0] delay_lane_e_20_sva;
  reg [4:0] delay_lane_e_10_sva;
  reg [4:0] delay_lane_e_21_sva;
  reg [4:0] delay_lane_e_9_sva;
  reg [4:0] delay_lane_e_22_sva;
  reg [4:0] delay_lane_e_8_sva;
  reg [4:0] delay_lane_e_23_sva;
  reg [4:0] delay_lane_e_7_sva;
  reg [4:0] delay_lane_e_24_sva;
  reg [4:0] delay_lane_e_6_sva;
  reg [4:0] delay_lane_e_25_sva;
  reg [4:0] delay_lane_e_5_sva;
  reg [4:0] delay_lane_e_26_sva;
  reg [4:0] delay_lane_e_4_sva;
  reg [4:0] delay_lane_e_27_sva;
  reg [4:0] delay_lane_e_3_sva;
  reg [4:0] delay_lane_e_28_sva;
  reg [4:0] delay_lane_e_2_sva;
  reg [4:0] delay_lane_e_29_sva;
  reg [4:0] delay_lane_e_1_sva;
  reg [4:0] delay_lane_e_30_sva;
  reg [4:0] delay_lane_e_0_sva;
  reg [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva;
  reg [1:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  reg MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm;
  reg MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm;
  reg MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm;
  reg MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm;
  reg MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm;
  reg MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm;
  reg MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm;
  reg MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm;
  reg MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm;
  reg MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm;
  reg MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm;
  reg MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  wire return_e_rsci_idat_mx0c1;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire [6:0] nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3;
  wire operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32;
  wire [10:0] MAC_ac_float_cctor_m_1_lpi_1_dfm_1;
  wire [3:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0;
  wire [3:0] result_m_1_lpi_1_dfm_1_10_7;
  reg [3:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0;
  reg [3:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_26_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_27_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_28_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_29_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_30_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_31_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_lpi_1_dfm_10_7;
  reg MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_10_7;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_12;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_14;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_13;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_15;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0;
  wire [6:0] operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2;
  reg [7:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc;
  wire or_482_ssc;
  wire [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4;
  wire MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4;
  wire [3:0] MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0;
  wire result_m_1_lpi_1_dfm_1_6;
  wire [1:0] result_m_1_lpi_1_dfm_1_5_4;
  wire [3:0] result_m_1_lpi_1_dfm_1_3_0;
  wire [5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt;
  wire [6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt;
  reg result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_6;
  reg [1:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_5_4;
  wire and_352_ssc;
  wire and_358_ssc;
  wire and_362_ssc;
  wire and_365_ssc;
  wire and_371_ssc;
  wire and_376_ssc;
  wire and_381_ssc;
  wire and_385_ssc;
  wire and_389_ssc;
  wire and_393_ssc;
  wire and_398_ssc;
  wire and_402_ssc;
  wire and_406_ssc;
  wire and_410_ssc;
  wire and_415_ssc;
  wire and_419_ssc;
  wire and_423_ssc;
  wire and_427_ssc;
  wire and_433_ssc;
  wire and_438_ssc;
  wire and_443_ssc;
  wire and_448_ssc;
  wire and_452_ssc;
  wire and_456_ssc;
  wire and_460_ssc;
  wire and_464_ssc;
  wire and_468_ssc;
  wire and_472_ssc;
  wire and_476_ssc;
  wire and_480_ssc;
  wire and_484_ssc;
  wire and_488_ssc;
  wire and_492_ssc;
  wire and_496_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse;
  wire MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse;
  wire nor_294_cse;
  wire nor_299_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse;
  wire or_385_rgt;
  wire and_517_rgt;
  wire and_76_rgt;
  wire or_379_rgt;
  wire and_512_rgt;
  wire nor_99_rgt;
  wire or_372_rgt;
  wire and_507_rgt;
  wire nor_100_rgt;
  wire or_369_rgt;
  wire and_503_rgt;
  wire nor_101_rgt;
  wire or_363_rgt;
  wire and_499_rgt;
  wire nor_102_rgt;
  wire or_292_rgt;
  wire and_343_rgt;
  wire nor_103_rgt;
  wire or_281_rgt;
  wire and_333_rgt;
  wire nor_104_rgt;
  wire or_275_rgt;
  wire and_329_rgt;
  wire and_85_rgt;
  wire or_268_rgt;
  wire and_325_rgt;
  wire and_87_rgt;
  wire or_260_rgt;
  wire and_321_rgt;
  wire and_89_rgt;
  wire or_253_rgt;
  wire and_317_rgt;
  wire and_91_rgt;
  wire or_246_rgt;
  wire and_313_rgt;
  wire and_92_rgt;
  wire or_239_rgt;
  wire and_309_rgt;
  wire and_93_rgt;
  wire or_231_rgt;
  wire and_305_rgt;
  wire and_94_rgt;
  wire or_287_rgt;
  wire and_339_rgt;
  wire nor_105_rgt;
  wire and_1120_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse;
  wire mux_127_itm;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_itm;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  wire MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1;
  reg MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0;
  reg [3:0] MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1;
  wire and_cse;
  wire and_901_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_m1c;

  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_31_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl;
  wire mux_291_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire or_381_nl;
  wire or_384_nl;
  wire or_383_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl;
  wire mux_282_nl;
  wire mux_281_nl;
  wire nor_181_nl;
  wire mux_280_nl;
  wire nand_nl;
  wire and_509_nl;
  wire mux_115_nl;
  wire mux_114_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl;
  wire mux_277_nl;
  wire mux_276_nl;
  wire mux_275_nl;
  wire mux_274_nl;
  wire or_371_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl;
  wire mux_271_nl;
  wire mux_270_nl;
  wire mux_269_nl;
  wire mux_268_nl;
  wire or_366_nl;
  wire mux_121_nl;
  wire mux_120_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire mux_263_nl;
  wire mux_262_nl;
  wire nor_172_nl;
  wire or_360_nl;
  wire mux_123_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl;
  wire mux_126_nl;
  wire mux_125_nl;
  wire mux_124_nl;
  wire or_164_nl;
  wire mux_224_nl;
  wire mux_223_nl;
  wire mux_222_nl;
  wire mux_221_nl;
  wire mux_220_nl;
  wire or_291_nl;
  wire mux_130_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire mux_207_nl;
  wire mux_206_nl;
  wire mux_205_nl;
  wire or_280_nl;
  wire or_279_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl;
  wire mux_201_nl;
  wire mux_200_nl;
  wire nor_159_nl;
  wire mux_199_nl;
  wire or_272_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl;
  wire mux_197_nl;
  wire nor_157_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire or_266_nl;
  wire or_264_nl;
  wire or_263_nl;
  wire mux_133_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl;
  wire mux_193_nl;
  wire nor_155_nl;
  wire mux_192_nl;
  wire mux_191_nl;
  wire or_258_nl;
  wire or_257_nl;
  wire mux_135_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl;
  wire MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl;
  wire mux_189_nl;
  wire nor_153_nl;
  wire mux_188_nl;
  wire mux_187_nl;
  wire or_251_nl;
  wire or_250_nl;
  wire mux_136_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl;
  wire MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl;
  wire mux_185_nl;
  wire nor_151_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire or_244_nl;
  wire or_243_nl;
  wire mux_137_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl;
  wire MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl;
  wire mux_181_nl;
  wire nor_149_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire or_237_nl;
  wire or_236_nl;
  wire mux_138_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl;
  wire MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl;
  wire mux_177_nl;
  wire mux_176_nl;
  wire nor_147_nl;
  wire mux_175_nl;
  wire or_228_nl;
  wire or_226_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl;
  wire MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl;
  wire MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl;
  wire MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl;
  wire mux_216_nl;
  wire mux_215_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire or_286_nl;
  wire mux_142_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl;
  wire mux_460_nl;
  wire mux_459_nl;
  wire mux_458_nl;
  wire mux_433_nl;
  wire mux_468_nl;
  wire mux_506_nl;
  wire and_900_nl;
  wire mux_429_nl;
  wire mux_428_nl;
  wire mux_465_nl;
  wire mux_507_nl;
  wire and_903_nl;
  wire mux_425_nl;
  wire mux_nl;
  wire and_890_nl;
  wire or_504_nl;
  wire or_nl;
  wire MAC_10_r_ac_float_else_and_nl;
  wire[4:0] MAC_10_r_ac_float_else_and_1_nl;
  wire mux_418_nl;
  wire mux_417_nl;
  wire mux_415_nl;
  wire mux_414_nl;
  wire mux_413_nl;
  wire mux_412_nl;
  wire mux_411_nl;
  wire mux_410_nl;
  wire mux_408_nl;
  wire mux_407_nl;
  wire mux_406_nl;
  wire mux_405_nl;
  wire mux_404_nl;
  wire mux_403_nl;
  wire mux_402_nl;
  wire mux_401_nl;
  wire mux_400_nl;
  wire mux_399_nl;
  wire mux_398_nl;
  wire mux_397_nl;
  wire mux_396_nl;
  wire mux_395_nl;
  wire mux_424_nl;
  wire mux_423_nl;
  wire mux_422_nl;
  wire mux_421_nl;
  wire and_889_nl;
  wire mux_505_nl;
  wire and_1148_nl;
  wire mux_504_nl;
  wire mux_503_nl;
  wire mux_502_nl;
  wire mux_501_nl;
  wire mux_500_nl;
  wire or_568_nl;
  wire mux_499_nl;
  wire mux_498_nl;
  wire mux_497_nl;
  wire mux_496_nl;
  wire mux_495_nl;
  wire mux_494_nl;
  wire mux_493_nl;
  wire mux_492_nl;
  wire mux_491_nl;
  wire mux_490_nl;
  wire mux_489_nl;
  wire mux_488_nl;
  wire mux_487_nl;
  wire mux_486_nl;
  wire mux_485_nl;
  wire mux_484_nl;
  wire mux_483_nl;
  wire mux_482_nl;
  wire mux_481_nl;
  wire mux_480_nl;
  wire mux_479_nl;
  wire mux_478_nl;
  wire mux_477_nl;
  wire mux_476_nl;
  wire mux_475_nl;
  wire mux_474_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire mux_367_nl;
  wire mux_366_nl;
  wire or_437_nl;
  wire and_665_nl;
  wire mux_371_nl;
  wire mux_370_nl;
  wire mux_149_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_nl;
  wire mux_364_nl;
  wire nor_209_nl;
  wire mux_363_nl;
  wire mux_362_nl;
  wire or_433_nl;
  wire and_661_nl;
  wire mux_365_nl;
  wire mux_151_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl;
  wire mux_360_nl;
  wire mux_359_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire or_428_nl;
  wire and_657_nl;
  wire mux_361_nl;
  wire mux_153_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_nl;
  wire mux_352_nl;
  wire mux_351_nl;
  wire mux_350_nl;
  wire nor_201_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire nor_204_nl;
  wire and_882_nl;
  wire and_653_nl;
  wire mux_353_nl;
  wire mux_155_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl;
  wire mux_346_nl;
  wire nor_198_nl;
  wire mux_345_nl;
  wire mux_344_nl;
  wire or_416_nl;
  wire and_649_nl;
  wire mux_347_nl;
  wire mux_156_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_nl;
  wire mux_342_nl;
  wire nor_195_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire or_412_nl;
  wire and_645_nl;
  wire mux_343_nl;
  wire mux_157_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl;
  wire mux_338_nl;
  wire nor_192_nl;
  wire mux_337_nl;
  wire mux_336_nl;
  wire or_408_nl;
  wire and_641_nl;
  wire mux_339_nl;
  wire mux_158_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_nl;
  wire mux_334_nl;
  wire nor_189_nl;
  wire mux_333_nl;
  wire mux_332_nl;
  wire or_404_nl;
  wire and_637_nl;
  wire mux_335_nl;
  wire mux_159_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_136_nl;
  wire mux_389_nl;
  wire mux_388_nl;
  wire or_478_nl;
  wire and_689_nl;
  wire mux_390_nl;
  wire mux_160_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl;
  wire mux_386_nl;
  wire nor_229_nl;
  wire mux_385_nl;
  wire or_471_nl;
  wire and_685_nl;
  wire mux_387_nl;
  wire mux_161_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl;
  wire mux_383_nl;
  wire nor_225_nl;
  wire mux_382_nl;
  wire or_464_nl;
  wire and_681_nl;
  wire mux_384_nl;
  wire mux_162_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_nl;
  wire mux_380_nl;
  wire nor_221_nl;
  wire mux_379_nl;
  wire or_457_nl;
  wire and_677_nl;
  wire mux_381_nl;
  wire mux_163_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_132_nl;
  wire mux_377_nl;
  wire mux_376_nl;
  wire mux_375_nl;
  wire or_450_nl;
  wire or_449_nl;
  wire and_673_nl;
  wire mux_378_nl;
  wire mux_164_nl;
  wire nor_114_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_16_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_30_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl;
  wire mux_373_nl;
  wire nor_216_nl;
  wire mux_372_nl;
  wire or_443_nl;
  wire and_669_nl;
  wire mux_374_nl;
  wire nor_93_nl;
  wire[2:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[3:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire MAC_3_r_ac_float_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_else_and_1_nl;
  wire mux_165_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_15_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_32_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl;
  wire mux_166_nl;
  wire mux_331_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[1:0] MAC_11_r_ac_float_else_and_nl;
  wire[3:0] MAC_11_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_12_r_ac_float_else_and_nl;
  wire[4:0] MAC_12_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_13_r_ac_float_else_and_nl;
  wire[4:0] MAC_13_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_14_r_ac_float_else_and_nl;
  wire[4:0] MAC_14_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_15_r_ac_float_else_and_nl;
  wire[4:0] MAC_15_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_16_r_ac_float_else_and_nl;
  wire[4:0] MAC_16_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_17_r_ac_float_else_and_nl;
  wire[4:0] MAC_17_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_2_r_ac_float_else_and_nl;
  wire[4:0] MAC_2_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_4_r_ac_float_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_5_r_ac_float_else_and_nl;
  wire[4:0] MAC_5_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_6_r_ac_float_else_and_nl;
  wire[4:0] MAC_6_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_7_r_ac_float_else_and_nl;
  wire[4:0] MAC_7_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_8_r_ac_float_else_and_nl;
  wire[4:0] MAC_8_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_9_r_ac_float_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_else_and_1_nl;
  wire MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire and_163_nl;
  wire and_166_nl;
  wire and_169_nl;
  wire MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire and_172_nl;
  wire and_175_nl;
  wire and_178_nl;
  wire MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_122_nl;
  wire and_185_nl;
  wire MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_123_nl;
  wire and_187_nl;
  wire MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire and_190_nl;
  wire and_193_nl;
  wire and_196_nl;
  wire MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_125_nl;
  wire and_198_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl;
  wire[3:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_126_nl;
  wire and_200_nl;
  wire MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_127_nl;
  wire and_202_nl;
  wire MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_128_nl;
  wire and_204_nl;
  wire MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_129_nl;
  wire and_206_nl;
  wire MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_130_nl;
  wire and_208_nl;
  wire MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_131_nl;
  wire and_210_nl;
  wire MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl;
  wire MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl;
  wire MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl;
  wire MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl;
  wire MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl;
  wire MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl;
  wire MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl;
  wire MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl;
  wire MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl;
  wire MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl;
  wire MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl;
  wire MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl;
  wire MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl;
  wire MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl;
  wire[3:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl;
  wire and_181_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[10:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_64_nl;
  wire[10:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[1:0] MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire MAC_18_r_ac_float_else_and_nl;
  wire[4:0] MAC_18_r_ac_float_else_and_1_nl;
  wire MAC_19_r_ac_float_else_and_nl;
  wire[4:0] MAC_19_r_ac_float_else_and_1_nl;
  wire MAC_20_r_ac_float_else_and_nl;
  wire[4:0] MAC_20_r_ac_float_else_and_1_nl;
  wire MAC_21_r_ac_float_else_and_nl;
  wire MAC_21_r_ac_float_else_and_1_nl;
  wire[3:0] MAC_21_r_ac_float_else_and_2_nl;
  wire MAC_22_r_ac_float_else_and_nl;
  wire[4:0] MAC_22_r_ac_float_else_and_1_nl;
  wire MAC_23_r_ac_float_else_and_nl;
  wire[4:0] MAC_23_r_ac_float_else_and_1_nl;
  wire MAC_24_r_ac_float_else_and_nl;
  wire[4:0] MAC_24_r_ac_float_else_and_1_nl;
  wire MAC_25_r_ac_float_else_and_nl;
  wire[4:0] MAC_25_r_ac_float_else_and_1_nl;
  wire MAC_26_r_ac_float_else_and_nl;
  wire[4:0] MAC_26_r_ac_float_else_and_1_nl;
  wire MAC_27_r_ac_float_else_and_nl;
  wire[4:0] MAC_27_r_ac_float_else_and_1_nl;
  wire MAC_28_r_ac_float_else_and_nl;
  wire[4:0] MAC_28_r_ac_float_else_and_1_nl;
  wire MAC_29_r_ac_float_else_and_nl;
  wire[4:0] MAC_29_r_ac_float_else_and_1_nl;
  wire MAC_30_r_ac_float_else_and_nl;
  wire[4:0] MAC_30_r_ac_float_else_and_1_nl;
  wire MAC_31_r_ac_float_else_and_nl;
  wire[4:0] MAC_31_r_ac_float_else_and_1_nl;
  wire MAC_1_r_ac_float_else_and_nl;
  wire[4:0] MAC_1_r_ac_float_else_and_1_nl;
  wire MAC_32_r_ac_float_else_and_nl;
  wire[4:0] MAC_32_r_ac_float_else_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl;
  wire[6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl;
  wire[6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl;
  wire[6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl;
  wire[6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl;
  wire[6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl;
  wire[6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl;
  wire[6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl;
  wire[6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl;
  wire[6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl;
  wire[6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl;
  wire[6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl;
  wire[6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl;
  wire[6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl;
  wire[6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl;
  wire[6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl;
  wire ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl;
  wire[5:0] MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_99_nl;
  wire[1:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_158_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_132_nl;
  wire[3:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_159_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_133_nl;
  wire[6:0] MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl;
  wire[7:0] nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl;
  wire[5:0] MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire mux_128_nl;
  wire mux_140_nl;
  wire or_189_nl;
  wire mux_171_nl;
  wire mux_170_nl;
  wire mux_169_nl;
  wire or_219_nl;
  wire mux_203_nl;
  wire mux_325_nl;
  wire mux_324_nl;
  wire mux_323_nl;
  wire mux_322_nl;
  wire or_392_nl;
  wire or_528_nl;
  wire or_540_nl;
  wire or_541_nl;
  wire or_542_nl;
  wire or_543_nl;
  wire or_544_nl;
  wire or_545_nl;
  wire or_546_nl;
  wire or_547_nl;
  wire or_548_nl;
  wire or_550_nl;
  wire mux_447_nl;
  wire mux_446_nl;
  wire or_549_nl;
  wire mux_450_nl;
  wire mux_449_nl;
  wire mux_436_nl;
  wire mux_453_nl;
  wire mux_452_nl;
  wire mux_470_nl;
  wire mux_435_nl;
  wire mux_509_nl;
  wire mux_456_nl;
  wire mux_455_nl;
  wire mux_432_nl;
  wire mux_508_nl;
  wire mux_434_nl;
  wire mux_427_nl;
  wire mux_471_nl;
  wire mux_230_nl;
  wire mux_229_nl;
  wire nor_30_nl;
  wire mux_261_nl;
  wire mux_260_nl;
  wire mux_259_nl;
  wire mux_258_nl;
  wire mux_257_nl;
  wire nor_171_nl;
  wire mux_256_nl;
  wire or_327_nl;
  wire or_326_nl;
  wire mux_255_nl;
  wire mux_254_nl;
  wire or_325_nl;
  wire or_324_nl;
  wire mux_253_nl;
  wire or_323_nl;
  wire or_322_nl;
  wire mux_252_nl;
  wire mux_251_nl;
  wire mux_250_nl;
  wire or_321_nl;
  wire or_320_nl;
  wire mux_249_nl;
  wire or_319_nl;
  wire or_318_nl;
  wire mux_248_nl;
  wire mux_247_nl;
  wire or_317_nl;
  wire or_316_nl;
  wire mux_246_nl;
  wire or_315_nl;
  wire or_314_nl;
  wire mux_245_nl;
  wire mux_244_nl;
  wire mux_243_nl;
  wire mux_242_nl;
  wire or_313_nl;
  wire or_312_nl;
  wire mux_241_nl;
  wire or_311_nl;
  wire or_310_nl;
  wire mux_240_nl;
  wire mux_239_nl;
  wire or_309_nl;
  wire or_308_nl;
  wire mux_238_nl;
  wire or_307_nl;
  wire or_306_nl;
  wire mux_237_nl;
  wire mux_236_nl;
  wire mux_235_nl;
  wire or_305_nl;
  wire or_304_nl;
  wire mux_234_nl;
  wire or_303_nl;
  wire or_302_nl;
  wire mux_233_nl;
  wire mux_232_nl;
  wire or_301_nl;
  wire or_300_nl;
  wire mux_231_nl;
  wire or_299_nl;
  wire or_298_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_32_nl;
  wire[4:0] and_905_nl;
  wire[4:0] mux1h_1_nl;
  wire[4:0] MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire and_696_nl;
  wire or_555_nl;
  wire mux_394_nl;
  wire nand_18_nl;
  wire or_489_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire mux_391_nl;
  wire or_502_nl;
  wire nor_237_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_96_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_97_nl;
  wire and_701_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_98_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_99_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_100_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_101_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_102_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_103_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_104_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_105_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_106_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_107_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_108_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_109_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_110_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_111_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_112_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_113_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_114_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_115_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_116_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_117_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_118_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_119_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_120_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_121_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_122_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_123_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_124_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_125_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_126_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_129_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_130_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_131_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_132_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_133_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_134_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_135_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_136_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_137_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_138_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_139_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_140_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_141_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_142_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_143_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_144_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_145_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_146_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_147_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_148_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_149_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_150_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_151_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_152_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_153_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_154_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_155_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_156_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_157_nl;
  wire not_995_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire and_898_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_128_nl;
  wire[3:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl;
  wire and_183_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_10_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_16_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl;
  wire[7:0] acc_nl;
  wire[8:0] nl_acc_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl;
  wire and_1151_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_158_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_159_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_160_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [12:0] nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl;
  wire [5:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2((MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_51_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_nl;
  wire [4:0] nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_51_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[4]), MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[3:0]), MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_51_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_54_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_nl;
  wire [4:0] nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_54_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[4]), MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[3:0]), MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_54_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_57_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_nl;
  wire [4:0] nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_57_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[4]), MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[3:0]), MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_57_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_60_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_nl;
  wire [4:0] nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_60_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg[4]), MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg[3:0]), MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_60_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_63_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_nl;
  wire [4:0] nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_63_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[4]), MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[3:0]), MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_63_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_66_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_nl;
  wire [4:0] nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_66_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[4]), MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[3:0]), MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_66_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_69_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_nl;
  wire [4:0] nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_69_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[4]), MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[3:0]), MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_69_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_72_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_nl;
  wire [4:0] nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_72_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[4]), MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[3:0]), MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_72_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_75_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_nl;
  wire [4:0] nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_75_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[4]), MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[3:0]), MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_75_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_78_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_nl;
  wire [4:0] nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_78_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[4]), MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[3:0]), MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_78_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_81_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_nl;
  wire [4:0] nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_81_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[4]), MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[3:0]), MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_81_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_84_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_nl;
  wire [4:0] nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_84_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[4]), MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[3:0]), MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_84_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_87_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_nl;
  wire [4:0] nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_87_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[4]), MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[3:0]), MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_87_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_90_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_nl;
  wire [4:0] nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_90_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[4]), MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[3:0]), MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_90_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_93_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_nl;
  wire [4:0] nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_93_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[4]), MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[3:0]), MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_93_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_nl};
  wire [11:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 , 1'b0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl;
  wire [5:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl
      , MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl;
  wire [5:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl;
  wire [5:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva;
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl
      , MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl;
  wire [5:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva;
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl;
  wire [5:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva;
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl
      , MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      , MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      , MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      , MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      , MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      , MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl;
  wire [5:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva;
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl
      , MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl;
  wire [5:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva;
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl
      , MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl;
  wire [5:0] nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva;
  assign nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl
      , MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , 1'b0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl;
  wire [5:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[1])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm};
  wire [4:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s;
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva};
  wire [12:0] nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_and_nl;
  wire [12:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_and_nl
      = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0]) & and_dcpl_59
      & (~ (fsm_output[5])) & (fsm_output[3]) & (~ (fsm_output[7])) & (fsm_output[0])
      & nor_294_cse;
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_and_nl};
  wire [12:0] nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd11)) input_m_rsci (
      .dat(input_m_rsc_dat),
      .idat(input_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd5)) input_e_rsci (
      .dat(input_e_rsc_dat),
      .idat(input_e_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd352)) taps_m_rsci (
      .dat(taps_m_rsc_dat),
      .idat(taps_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd160)) taps_e_rsci (
      .dat(taps_e_rsc_dat),
      .idat(taps_e_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd5),
  .width(32'sd11)) return_m_rsci (
      .idat(return_m_rsci_idat),
      .dat(return_m_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd6),
  .width(32'sd5)) return_e_rsci (
      .idat(return_e_rsci_idat),
      .dat(return_e_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_m_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(input_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_e_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(input_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_m_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(taps_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_e_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(taps_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_m_triosy_obj (
      .ld(reg_return_e_triosy_obj_ld_cse),
      .lz(return_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_e_triosy_obj (
      .ld(reg_return_e_triosy_obj_ld_cse),
      .lz(return_e_triosy_lz)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1),
      .z(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva),
      .s(nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1),
      .z(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva),
      .s(nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1),
      .z(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva),
      .s(nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1),
      .z(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva),
      .s(nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1),
      .z(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva),
      .s(nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1),
      .z(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva),
      .s(nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1),
      .z(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva),
      .s(nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1),
      .z(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva),
      .s(nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1),
      .z(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva),
      .s(nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1),
      .z(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva),
      .s(nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1),
      .z(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva),
      .s(nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1),
      .z(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva),
      .s(nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1),
      .z(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva),
      .s(nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1),
      .z(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva),
      .s(nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1),
      .z(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[11:0]),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva),
      .s(nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm),
      .z(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_12),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_14)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s[4:0]),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  leading_sign_13_1_1_0  MAC_10_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_13),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_15)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_2)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_4)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_5)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_6)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_7)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_8)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_9)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_10)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_11)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_12)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_13)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0),
      .z(z_out_14)
    );
  fir_core_wait_dp fir_core_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse = and_dcpl_64
      | and_dcpl_67;
  assign or_138_cse = (fsm_output[2:1]!=2'b00);
  assign nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_30_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[154:150]);
  assign MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_381_nl = (fsm_output[3]) | (~ or_tmp_62);
  assign mux_289_nl = MUX_s_1_2_2(mux_tmp_284, or_381_nl, fsm_output[2]);
  assign or_384_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[5:4]!=2'b00);
  assign mux_290_nl = MUX_s_1_2_2(mux_tmp_285, mux_289_nl, or_384_nl);
  assign or_383_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[6]);
  assign mux_291_nl = MUX_s_1_2_2(mux_290_nl, mux_tmp_285, or_383_nl);
  assign or_385_rgt = mux_291_nl | or_dcpl_170;
  assign and_517_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm))
      & and_dcpl_93 & and_dcpl_343;
  assign and_76_rgt = (~((~(or_138_cse ^ (fsm_output[3]))) | (fsm_output[7]))) &
      (fsm_output[6:4]==3'b000);
  assign nor_179_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[4]));
  assign nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_24_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[124:120]);
  assign MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nand_nl = ~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
      | (~ (fsm_output[0])))) & (~(nor_179_cse | (fsm_output[6]))));
  assign mux_280_nl = MUX_s_1_2_2((fsm_output[6]), nand_nl, fsm_output[1]);
  assign nor_181_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_280_nl);
  assign and_509_nl = (fsm_output[4]) & or_138_cse & (fsm_output[6]);
  assign mux_281_nl = MUX_s_1_2_2(nor_181_nl, and_509_nl, fsm_output[3]);
  assign mux_282_nl = MUX_s_1_2_2(mux_281_nl, (fsm_output[6]), fsm_output[5]);
  assign or_379_rgt = mux_282_nl | (fsm_output[7]);
  assign and_512_rgt = (nor_179_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_114_nl = MUX_s_1_2_2((~ or_tmp_92), mux_tmp_110, fsm_output[4]);
  assign mux_115_nl = MUX_s_1_2_2(mux_114_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_99_rgt = ~(mux_115_nl | (fsm_output[7]));
  assign nor_177_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5);
  assign nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_23_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[119:115]);
  assign MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_371_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[4]);
  assign mux_274_nl = MUX_s_1_2_2(or_tmp_92, or_tmp_204, or_371_nl);
  assign mux_275_nl = MUX_s_1_2_2(mux_274_nl, or_tmp_92, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6);
  assign mux_276_nl = MUX_s_1_2_2((~ mux_275_nl), mux_tmp_113, fsm_output[4]);
  assign mux_277_nl = MUX_s_1_2_2(mux_276_nl, (fsm_output[6]), fsm_output[5]);
  assign or_372_rgt = mux_277_nl | (fsm_output[7]);
  assign and_507_rgt = (nor_177_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_117_nl = MUX_s_1_2_2((~ or_tmp_92), mux_tmp_113, fsm_output[4]);
  assign mux_118_nl = MUX_s_1_2_2(mux_117_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_100_rgt = ~(mux_118_nl | (fsm_output[7]));
  assign nor_175_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5);
  assign or_92_cse = (fsm_output[3:2]!=2'b00);
  assign nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_22_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[114:110]);
  assign MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_366_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[4]);
  assign mux_268_nl = MUX_s_1_2_2(or_tmp_92, or_tmp_204, or_366_nl);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, or_tmp_92, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6);
  assign mux_270_nl = MUX_s_1_2_2((~ mux_269_nl), mux_tmp_116, fsm_output[4]);
  assign mux_271_nl = MUX_s_1_2_2(mux_270_nl, (fsm_output[6]), fsm_output[5]);
  assign or_369_rgt = mux_271_nl | (fsm_output[7]);
  assign and_503_rgt = (nor_175_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_120_nl = MUX_s_1_2_2((~ or_tmp_92), mux_tmp_116, fsm_output[4]);
  assign mux_121_nl = MUX_s_1_2_2(mux_120_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_101_rgt = ~(mux_121_nl | (fsm_output[7]));
  assign or_359_cse = (fsm_output[5:4]!=2'b00);
  assign nor_173_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5);
  assign and_867_cse = (fsm_output[3]) & (fsm_output[1]) & (fsm_output[6]);
  assign nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_21_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[109:105]);
  assign MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nor_172_nl = ~((fsm_output[6]) | (fsm_output[3]) | (~ or_tmp_100));
  assign mux_262_nl = MUX_s_1_2_2(nor_172_nl, and_867_cse, fsm_output[2]);
  assign or_360_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[4]);
  assign mux_263_nl = MUX_s_1_2_2(mux_tmp_119, mux_262_nl, or_360_nl);
  assign mux_264_nl = MUX_s_1_2_2(mux_263_nl, mux_tmp_119, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, (fsm_output[6]), or_359_cse);
  assign or_363_rgt = mux_265_nl | (fsm_output[7]);
  assign and_499_rgt = (nor_173_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_123_nl = MUX_s_1_2_2(mux_tmp_119, (fsm_output[6]), or_359_cse);
  assign nor_102_rgt = ~(mux_123_nl | (fsm_output[7]));
  assign or_165_cse = (fsm_output[6]) | (fsm_output[3]);
  assign nor_169_cse = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1!=2'b00));
  assign nor_66_cse = ~((fsm_output[0]) | (fsm_output[7]));
  assign and_880_cse = (fsm_output[1:0]==2'b11);
  assign nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_20_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[104:100]);
  assign MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_125_nl = MUX_s_1_2_2(or_tmp_100, or_tmp_96, or_165_cse);
  assign or_164_nl = and_880_cse | (fsm_output[7]);
  assign mux_124_nl = MUX_s_1_2_2(or_164_nl, or_tmp_96, or_165_cse);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, mux_124_nl, fsm_output[2]);
  assign mux_127_itm = MUX_s_1_2_2(mux_126_nl, or_tmp_96, or_359_cse);
  assign nor_166_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5);
  assign nor_61_cse = ~((fsm_output[3]) | (fsm_output[6]));
  assign nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_19_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[99:95]);
  assign MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_220_nl = MUX_s_1_2_2((~ or_tmp_128), nor_tmp_24, fsm_output[6]);
  assign mux_221_nl = MUX_s_1_2_2(mux_220_nl, nor_tmp_12, fsm_output[2]);
  assign or_291_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[4]);
  assign mux_222_nl = MUX_s_1_2_2(mux_tmp_126, mux_221_nl, or_291_nl);
  assign mux_223_nl = MUX_s_1_2_2(mux_222_nl, mux_tmp_126, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6);
  assign mux_224_nl = MUX_s_1_2_2(mux_223_nl, (fsm_output[6]), or_359_cse);
  assign or_292_rgt = mux_224_nl | (fsm_output[7]);
  assign and_343_rgt = (nor_166_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_130_nl = MUX_s_1_2_2(mux_tmp_126, (fsm_output[6]), or_359_cse);
  assign nor_103_rgt = ~(mux_130_nl | (fsm_output[7]));
  assign nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_18_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[94:90]);
  assign MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_205_nl = MUX_s_1_2_2((~ or_tmp_128), or_tmp_25, fsm_output[6]);
  assign mux_206_nl = MUX_s_1_2_2(mux_205_nl, (fsm_output[6]), fsm_output[2]);
  assign or_280_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[5:4]!=2'b00);
  assign mux_207_nl = MUX_s_1_2_2(mux_tmp_201, mux_206_nl, or_280_nl);
  assign or_279_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[6]);
  assign mux_208_nl = MUX_s_1_2_2(mux_207_nl, mux_tmp_201, or_279_nl);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, (fsm_output[6]), or_359_cse);
  assign or_281_rgt = mux_209_nl | (fsm_output[7]);
  assign and_333_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign nor_104_rgt = ~((~((or_dcpl_66 | or_359_cse) ^ (fsm_output[6]))) | (fsm_output[7]));
  assign nor_160_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[5:4]!=2'b00));
  assign nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_17_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[89:85]);
  assign MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_199_nl = MUX_s_1_2_2(or_tmp_25, or_tmp_128, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm);
  assign nor_159_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_199_nl);
  assign mux_200_nl = MUX_s_1_2_2(nor_159_nl, nor_tmp_9, fsm_output[5]);
  assign or_272_nl = nor_160_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[6]);
  assign mux_201_nl = MUX_s_1_2_2(mux_200_nl, mux_tmp_128, or_272_nl);
  assign or_275_rgt = mux_201_nl | or_dcpl_100;
  assign and_329_rgt = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[6])
      | nor_160_cse) & and_dcpl_93 & and_dcpl_290;
  assign and_85_rgt = (~ mux_tmp_128) & and_dcpl_1;
  assign nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_16_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[84:80]);
  assign MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_266_nl = (fsm_output[3:2]!=2'b00) | (~ or_tmp_100);
  assign or_264_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[5:4]!=2'b00);
  assign mux_195_nl = MUX_s_1_2_2(or_dcpl_66, or_266_nl, or_264_nl);
  assign or_263_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[6]);
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, or_dcpl_66, or_263_nl);
  assign nor_157_nl = ~((fsm_output[4]) | mux_196_nl);
  assign mux_197_nl = MUX_s_1_2_2(nor_157_nl, and_tmp_6, fsm_output[5]);
  assign or_268_rgt = mux_197_nl | or_dcpl_100;
  assign and_325_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign mux_133_nl = MUX_s_1_2_2(or_tmp_102, (~ and_tmp_6), fsm_output[5]);
  assign and_87_rgt = mux_133_nl & and_dcpl_1;
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_15_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_258_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[5:4]!=2'b00);
  assign mux_191_nl = MUX_s_1_2_2(or_tmp_25, or_tmp_128, or_258_nl);
  assign or_257_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[6]);
  assign mux_192_nl = MUX_s_1_2_2(mux_191_nl, or_tmp_25, or_257_nl);
  assign nor_155_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_192_nl);
  assign mux_193_nl = MUX_s_1_2_2(nor_155_nl, and_tmp_7, fsm_output[5]);
  assign or_260_rgt = mux_193_nl | or_dcpl_100;
  assign and_321_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign mux_135_nl = MUX_s_1_2_2(or_tmp_102, (~ and_tmp_7), fsm_output[5]);
  assign and_89_rgt = mux_135_nl & and_dcpl_1;
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_14_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_251_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[5:4]!=2'b00);
  assign mux_187_nl = MUX_s_1_2_2(or_tmp_25, or_tmp_128, or_251_nl);
  assign or_250_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[6]);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, or_tmp_25, or_250_nl);
  assign nor_153_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_188_nl);
  assign mux_189_nl = MUX_s_1_2_2(nor_153_nl, and_tmp_8, fsm_output[5]);
  assign or_253_rgt = mux_189_nl | or_dcpl_100;
  assign and_317_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign mux_136_nl = MUX_s_1_2_2(or_tmp_102, (~ and_tmp_8), fsm_output[5]);
  assign and_91_rgt = mux_136_nl & and_dcpl_1;
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_13_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_244_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[5:4]!=2'b00);
  assign mux_183_nl = MUX_s_1_2_2(or_tmp_25, or_tmp_128, or_244_nl);
  assign or_243_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[6]);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, or_tmp_25, or_243_nl);
  assign nor_151_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_184_nl);
  assign mux_185_nl = MUX_s_1_2_2(nor_151_nl, or_tmp_17, fsm_output[5]);
  assign or_246_rgt = mux_185_nl | or_dcpl_100;
  assign and_313_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign mux_137_nl = MUX_s_1_2_2(or_tmp_102, (~ or_tmp_17), fsm_output[5]);
  assign and_92_rgt = mux_137_nl & and_dcpl_1;
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_12_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_237_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[5:4]!=2'b00);
  assign mux_179_nl = MUX_s_1_2_2(or_tmp_25, or_tmp_128, or_237_nl);
  assign or_236_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[6]);
  assign mux_180_nl = MUX_s_1_2_2(mux_179_nl, or_tmp_25, or_236_nl);
  assign nor_149_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_180_nl);
  assign mux_181_nl = MUX_s_1_2_2(nor_149_nl, or_tmp_104, fsm_output[5]);
  assign or_239_rgt = mux_181_nl | or_dcpl_100;
  assign and_309_rgt = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm))
      & and_dcpl_93 & and_dcpl_290;
  assign mux_138_nl = MUX_s_1_2_2(or_tmp_102, (~ or_tmp_104), fsm_output[5]);
  assign and_93_rgt = mux_138_nl & and_dcpl_1;
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_11_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_228_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[6]);
  assign mux_175_nl = MUX_s_1_2_2(or_tmp_128, or_tmp_25, or_228_nl);
  assign nor_147_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_175_nl);
  assign mux_176_nl = MUX_s_1_2_2(nor_147_nl, or_tmp_105, fsm_output[5]);
  assign or_226_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[5:4]!=2'b00);
  assign mux_177_nl = MUX_s_1_2_2(mux_tmp_136, mux_176_nl, or_226_nl);
  assign or_231_rgt = mux_177_nl | or_dcpl_100;
  assign and_305_rgt = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[5:4]!=2'b00))))
      & and_dcpl_93 & and_dcpl_290;
  assign and_94_rgt = (~ mux_tmp_136) & and_dcpl_1;
  assign nor_164_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5);
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(input_e_rsci_idat)
      + conv_s2s_5_6(taps_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_212_nl = MUX_s_1_2_2((~ or_tmp_128), (fsm_output[3]), fsm_output[6]);
  assign mux_213_nl = MUX_s_1_2_2(mux_212_nl, and_tmp_3, fsm_output[2]);
  assign or_286_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[4]);
  assign mux_214_nl = MUX_s_1_2_2(mux_tmp_138, mux_213_nl, or_286_nl);
  assign mux_215_nl = MUX_s_1_2_2(mux_214_nl, mux_tmp_138, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6);
  assign mux_216_nl = MUX_s_1_2_2(mux_215_nl, (fsm_output[6]), or_359_cse);
  assign or_287_rgt = mux_216_nl | (fsm_output[7]);
  assign and_339_rgt = (nor_164_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6)
      & and_dcpl_98 & and_dcpl_324;
  assign mux_142_nl = MUX_s_1_2_2(mux_tmp_138, (fsm_output[6]), or_359_cse);
  assign nor_105_rgt = ~(mux_142_nl | (fsm_output[7]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
      = (~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_91;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse
      = MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_91;
  assign or_183_cse = (fsm_output[6:2]!=5'b00000);
  assign and_698_m1c = and_dcpl_66 & and_dcpl_90;
  assign and_703_m1c = and_dcpl_688 & and_dcpl_60;
  assign and_704_m1c = and_dcpl_688 & and_dcpl_90;
  assign and_705_m1c = and_dcpl_66 & and_dcpl_514;
  assign and_706_m1c = and_dcpl_66 & and_dcpl_518;
  assign and_707_m1c = and_dcpl_688 & and_dcpl_514;
  assign and_708_m1c = and_dcpl_688 & and_dcpl_518;
  assign and_709_m1c = and_dcpl_66 & and_dcpl_529;
  assign and_710_m1c = and_dcpl_66 & and_dcpl_533;
  assign and_711_m1c = and_dcpl_688 & and_dcpl_529;
  assign and_712_m1c = and_dcpl_688 & and_dcpl_533;
  assign and_713_m1c = and_dcpl_66 & and_dcpl_543;
  assign and_714_m1c = and_dcpl_66 & and_dcpl_547;
  assign and_715_m1c = and_dcpl_688 & and_dcpl_543;
  assign and_716_m1c = and_dcpl_688 & and_dcpl_547;
  assign and_717_m1c = and_dcpl_66 & and_dcpl_558;
  assign and_718_m1c = and_dcpl_66 & and_dcpl_570;
  assign and_719_m1c = and_dcpl_688 & and_dcpl_558;
  assign and_720_m1c = and_dcpl_688 & and_dcpl_570;
  assign and_721_m1c = and_dcpl_66 & and_dcpl_574;
  assign and_722_m1c = and_dcpl_66 & and_dcpl_578;
  assign and_723_m1c = and_dcpl_688 & and_dcpl_574;
  assign and_724_m1c = and_dcpl_688 & and_dcpl_578;
  assign and_725_m1c = and_dcpl_66 & and_dcpl_589;
  assign and_726_m1c = and_dcpl_66 & and_dcpl_593;
  assign and_727_m1c = and_dcpl_688 & and_dcpl_589;
  assign and_728_m1c = and_dcpl_688 & and_dcpl_593;
  assign and_729_m1c = and_dcpl_66 & and_dcpl_609;
  assign and_730_m1c = and_dcpl_66 & and_dcpl_613;
  assign and_731_m1c = and_dcpl_688 & and_dcpl_609;
  assign and_732_m1c = and_dcpl_688 & and_dcpl_613;
  assign and_899_cse = and_dcpl_558 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  assign and_902_cse = and_dcpl_558 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva;
  assign and_cse = and_dcpl_90 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm;
  assign and_901_cse = and_dcpl_90 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  assign mux_506_nl = MUX_s_1_2_2(mux_tmp_427, or_tmp_270, and_cse);
  assign mux_468_nl = MUX_s_1_2_2(mux_506_nl, or_tmp_270, and_899_cse);
  assign and_900_nl = and_dcpl_578 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm;
  assign mux_433_nl = MUX_s_1_2_2(mux_468_nl, or_tmp_270, and_900_nl);
  assign mux_458_nl = MUX_s_1_2_2(mux_tmp_454, mux_433_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign mux_507_nl = MUX_s_1_2_2(or_tmp_283, or_tmp_270, and_901_cse);
  assign mux_465_nl = MUX_s_1_2_2(mux_507_nl, or_tmp_270, and_902_cse);
  assign and_903_nl = and_dcpl_578 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva;
  assign mux_428_nl = MUX_s_1_2_2(mux_465_nl, or_tmp_270, and_903_nl);
  assign mux_429_nl = MUX_s_1_2_2(mux_428_nl, or_tmp_270, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign mux_459_nl = MUX_s_1_2_2(mux_458_nl, mux_429_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm);
  assign mux_460_nl = MUX_s_1_2_2(mux_tmp_454, mux_459_nl, and_dcpl_593);
  assign and_890_nl = and_dcpl_66 & (and_dcpl_514 | and_dcpl_518 | and_dcpl_529 |
      and_dcpl_547 | and_dcpl_533 | and_dcpl_543 | and_dcpl_570 | and_dcpl_574 |
      and_dcpl_589 | and_dcpl_609 | and_dcpl_613);
  assign or_504_nl = and_dcpl_60 | and_dcpl_514 | and_dcpl_518 | and_dcpl_529 | and_dcpl_547
      | and_dcpl_533 | and_dcpl_543 | and_dcpl_570 | and_dcpl_574 | and_dcpl_589
      | and_dcpl_609 | and_dcpl_613;
  assign mux_nl = MUX_s_1_2_2(and_890_nl, or_504_nl, and_dcpl_688);
  assign or_nl = and_dcpl_593 | and_dcpl_578 | and_dcpl_558 | and_dcpl_90;
  assign mux_425_nl = MUX_s_1_2_2(mux_nl, or_tmp_270, or_nl);
  assign mux_461_tmp = MUX_s_1_2_2(mux_460_nl, mux_425_nl, MAC_3_result_operator_result_operator_nor_tmp);
  assign MAC_10_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      & MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_10_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2,
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm
      = conv_s2s_6_7({MAC_10_r_ac_float_else_and_nl , MAC_10_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6:0];
  assign mux_420_cse = MUX_s_1_2_2((MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_418_nl = MUX_s_1_2_2((MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_417_nl = MUX_s_1_2_2((MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_419_cse = MUX_s_1_2_2(mux_418_nl, mux_417_nl, fsm_output[6]);
  assign mux_414_nl = MUX_s_1_2_2((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_413_nl = MUX_s_1_2_2((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_415_nl = MUX_s_1_2_2(mux_414_nl, mux_413_nl, fsm_output[6]);
  assign mux_411_nl = MUX_s_1_2_2((MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_410_nl = MUX_s_1_2_2((MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_412_nl = MUX_s_1_2_2(mux_411_nl, mux_410_nl, fsm_output[6]);
  assign mux_416_cse = MUX_s_1_2_2(mux_415_nl, mux_412_nl, fsm_output[2]);
  assign mux_406_nl = MUX_s_1_2_2((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_405_nl = MUX_s_1_2_2((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_407_nl = MUX_s_1_2_2(mux_406_nl, mux_405_nl, fsm_output[6]);
  assign mux_403_nl = MUX_s_1_2_2((MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_402_nl = MUX_s_1_2_2((MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_404_nl = MUX_s_1_2_2(mux_403_nl, mux_402_nl, fsm_output[6]);
  assign mux_408_nl = MUX_s_1_2_2(mux_407_nl, mux_404_nl, fsm_output[2]);
  assign mux_399_nl = MUX_s_1_2_2((MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_398_nl = MUX_s_1_2_2((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_400_nl = MUX_s_1_2_2(mux_399_nl, mux_398_nl, fsm_output[6]);
  assign mux_396_nl = MUX_s_1_2_2((MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_395_nl = MUX_s_1_2_2((MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[3]);
  assign mux_397_nl = MUX_s_1_2_2(mux_396_nl, mux_395_nl, fsm_output[6]);
  assign mux_401_nl = MUX_s_1_2_2(mux_400_nl, mux_397_nl, fsm_output[2]);
  assign mux_409_cse = MUX_s_1_2_2(mux_408_nl, mux_401_nl, fsm_output[5]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_ssc = and_dcpl_64 | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1
      | and_dcpl_103 | and_dcpl_99;
  assign and_889_nl = (fsm_output[3]) & (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_421_nl = MUX_s_1_2_2(and_889_nl, mux_420_cse, fsm_output[6]);
  assign mux_422_nl = MUX_s_1_2_2(mux_421_nl, mux_419_cse, fsm_output[2]);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, mux_416_cse, fsm_output[5]);
  assign mux_424_nl = MUX_s_1_2_2(mux_423_nl, mux_409_cse, fsm_output[4]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse = mux_424_nl & and_dcpl_135;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_90;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse = and_dcpl_135 & (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_60 & and_dcpl_103;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_90;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_514;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_518;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse = and_dcpl_524 & (~((fsm_output[2])
      | (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_365;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_518;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_529;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_533;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_529;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_533;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_543;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_547;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_543;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_547;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_558;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse = and_dcpl_100 & and_dcpl_570;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse = and_dcpl_564 & and_dcpl_341
      & (~((fsm_output[5]) | (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_558;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_570;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_574;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_578;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_574;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse = and_dcpl_587 & (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & (fsm_output[2]) & and_dcpl_365;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_589;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse = and_dcpl_135 & (~((fsm_output[3])
      | (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_593;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse = and_dcpl_587 & (~((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[2]))) & and_dcpl_382;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse = and_dcpl_587 & (fsm_output[2])
      & (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_382;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse = and_dcpl_564 & (~((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[2]))) & and_dcpl_399;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse = and_dcpl_564 & (fsm_output[2])
      & (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_399;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_609;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse = and_dcpl_135 & (fsm_output[3])
      & (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_613;
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse = and_dcpl_148 | (and_dcpl_724
      & and_dcpl_60);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse = (and_dcpl_724 & and_dcpl_90)
      | (and_dcpl_724 & and_dcpl_613);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse = (and_dcpl_100 & and_dcpl_514)
      | (and_dcpl_724 & and_dcpl_609);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse = (and_dcpl_100 & and_dcpl_518)
      | (and_dcpl_100 & and_dcpl_613);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse = (and_dcpl_724 & and_dcpl_514)
      | (and_dcpl_100 & and_dcpl_609);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse = (and_dcpl_724 & and_dcpl_518)
      | (and_dcpl_724 & and_dcpl_593);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse = (and_dcpl_100 & and_dcpl_529)
      | (and_dcpl_724 & and_dcpl_589);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse = (and_dcpl_100 & and_dcpl_533)
      | (and_dcpl_100 & and_dcpl_593);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse = (and_dcpl_724 & and_dcpl_529)
      | (and_dcpl_100 & and_dcpl_589);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse = (and_dcpl_724 & and_dcpl_533)
      | (and_dcpl_724 & and_dcpl_578);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse = (and_dcpl_100 & and_dcpl_543)
      | (and_dcpl_724 & and_dcpl_574);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse = (and_dcpl_100 & and_dcpl_547)
      | (and_dcpl_100 & and_dcpl_578);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse = (and_dcpl_724 & and_dcpl_543)
      | (and_dcpl_100 & and_dcpl_574);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse = (and_dcpl_724 & and_dcpl_547)
      | (and_dcpl_724 & and_dcpl_570);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse = (and_dcpl_100 & and_dcpl_558)
      | (and_dcpl_724 & and_dcpl_558);
  assign or_553_tmp = ((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]))
      & (~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_67 & ((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm)
      | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva[21]) | (~ MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1]))
      & and_dcpl_95);
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg)}) +
      7'b0000001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_ssc = ~(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva[21]))
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_146_nl = MUX_s_1_2_2((~ or_tmp_110), nor_tmp_27, fsm_output[4]);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, (fsm_output[6]), fsm_output[5]);
  assign nor_106_ssc = ~(mux_147_nl | (fsm_output[7]));
  assign nor_212_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5);
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg)}) +
      7'b0000001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_ssc = ~(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva[21]))
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_149_nl = MUX_s_1_2_2(not_tmp_131, mux_tmp_145, fsm_output[5]);
  assign nor_107_ssc = ~(mux_149_nl | (fsm_output[7]));
  assign nor_210_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5);
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg)}) +
      7'b0000001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_ssc = ~(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva[21]))
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_151_nl = MUX_s_1_2_2(not_tmp_131, mux_tmp_147, fsm_output[5]);
  assign nor_108_ssc = ~(mux_151_nl | (fsm_output[7]));
  assign nor_207_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5);
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg)}) +
      7'b0000001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_ssc = ~(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva[21]))
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_153_nl = MUX_s_1_2_2(not_tmp_131, mux_tmp_149, fsm_output[5]);
  assign nor_109_ssc = ~(mux_153_nl | (fsm_output[7]));
  assign nor_202_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[4]));
  assign nor_203_cse = ~((fsm_output[6:5]!=2'b00));
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg)}) +
      7'b0000001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_ssc = ~(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva[21]))
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_155_nl = MUX_s_1_2_2(not_tmp_131, mux_tmp_151, fsm_output[5]);
  assign nor_110_ssc = ~(mux_155_nl | (fsm_output[7]));
  assign nor_199_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5);
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg)}) +
      7'b0000001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_ssc = ~(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva[21]))
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_156_nl = MUX_s_1_2_2(not_tmp_131, and_tmp_9, fsm_output[5]);
  assign nor_111_ssc = ~(mux_156_nl | (fsm_output[7]));
  assign nor_196_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5);
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg)}) + 7'b0000001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_ssc = ~(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva[21]))
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_157_nl = MUX_s_1_2_2(not_tmp_131, and_tmp_10, fsm_output[5]);
  assign nor_112_ssc = ~(mux_157_nl | (fsm_output[7]));
  assign nor_193_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5);
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg)}) + 7'b0000001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1);
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_ssc = ~(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva[21]))
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_158_nl = MUX_s_1_2_2(not_tmp_131, and_tmp_11, fsm_output[5]);
  assign nor_113_ssc = ~(mux_158_nl | (fsm_output[7]));
  assign nor_190_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5);
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg)}) + 7'b0000001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1);
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_ssc = ~(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva[21]))
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_159_nl = MUX_s_1_2_2(or_tmp_114, (~ nor_tmp_24), fsm_output[2]);
  assign and_129_ssc = mux_159_nl & and_dcpl_1 & and_dcpl_36;
  assign nor_231_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[5:4]!=2'b00));
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg)}) + 7'b0000001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1);
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_ssc = ~(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva[21]))
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_160_nl = MUX_s_1_2_2(or_tmp_116, (~ or_dcpl_66), fsm_output[4]);
  assign and_131_ssc = mux_160_nl & and_dcpl_118;
  assign nor_227_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[5:4]!=2'b00));
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg)}) + 7'b0000001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1);
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_ssc = ~(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva[21]))
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_161_nl = MUX_s_1_2_2(or_tmp_116, (~ mux_tmp_131), fsm_output[4]);
  assign and_132_ssc = mux_161_nl & and_dcpl_118;
  assign nor_223_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[5:4]!=2'b00));
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg)}) + 7'b0000001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1);
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_ssc = ~(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva[21]))
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_162_nl = MUX_s_1_2_2(or_tmp_116, (~ mux_tmp_129), fsm_output[4]);
  assign and_133_ssc = mux_162_nl & and_dcpl_118;
  assign nor_219_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[5:4]!=2'b00));
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg)}) + 7'b0000001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1);
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_ssc = ~(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva[21]))
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_163_nl = MUX_s_1_2_2(or_tmp_116, (~ and_861_cse), fsm_output[4]);
  assign and_134_ssc = mux_163_nl & and_dcpl_118;
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg)}) + 7'b0000001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1);
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_ssc = ~(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva[21]))
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign nor_114_nl = ~((fsm_output[4:2]!=3'b000) | and_880_cse);
  assign mux_164_nl = MUX_s_1_2_2(nor_114_nl, or_tmp_102, fsm_output[5]);
  assign and_135_ssc = (~ mux_164_nl) & and_dcpl_1;
  assign nor_214_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[5:4]!=2'b00));
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg)}) + 7'b0000001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1);
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_ssc = ~(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva[21]))
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign nor_187_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4])
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[0]));
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc = and_dcpl_129 | and_dcpl_95
      | and_dcpl_132;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse = and_dcpl_129 | and_dcpl_95;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse = ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse
      & (~ and_dcpl_67);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse
      = and_dcpl_67 | and_dcpl_95;
  assign MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse = ~((z_out_17!=11'b00000000000));
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc = and_dcpl_67
      | and_dcpl_91 | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_64_nl = ~ MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      = MUX_v_11_2_2(11'b00000000000, MAC_ac_float_cctor_m_1_lpi_1_dfm_1, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_64_nl);
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      = MUX_v_11_2_2(11'b00000000000, MAC_ac_float_cctor_m_1_lpi_1_dfm_1, MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = conv_s2u_11_12(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl)
      + conv_s2u_11_12(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl);
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[11:1])
      + conv_s2u_11_12({result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_10_7
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_6 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_5_4
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0});
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0 = $signed((input_m_rsci_idat))
      * $signed((taps_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0 = $signed(delay_lane_m_17_sva)
      * $signed((taps_m_rsci_idat[197:187]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0 = $signed(delay_lane_m_18_sva)
      * $signed((taps_m_rsci_idat[208:198]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0 = $signed(delay_lane_m_19_sva)
      * $signed((taps_m_rsci_idat[219:209]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0 = $signed(delay_lane_m_20_sva)
      * $signed((taps_m_rsci_idat[230:220]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0 = $signed(delay_lane_m_21_sva)
      * $signed((taps_m_rsci_idat[241:231]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0 = $signed(delay_lane_m_22_sva)
      * $signed((taps_m_rsci_idat[252:242]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0 = $signed(delay_lane_m_23_sva)
      * $signed((taps_m_rsci_idat[263:253]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0 = $signed(delay_lane_m_24_sva)
      * $signed((taps_m_rsci_idat[274:264]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0 = $signed(delay_lane_m_25_sva)
      * $signed((taps_m_rsci_idat[285:275]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0 = $signed(delay_lane_m_26_sva)
      * $signed((taps_m_rsci_idat[296:286]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0 = $signed(delay_lane_m_27_sva)
      * $signed((taps_m_rsci_idat[307:297]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0 = $signed(delay_lane_m_28_sva)
      * $signed((taps_m_rsci_idat[318:308]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0 = $signed(delay_lane_m_29_sva)
      * $signed((taps_m_rsci_idat[329:319]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0 = $signed(delay_lane_m_30_sva)
      * $signed((taps_m_rsci_idat[340:330]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0 = $signed(({MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7
      , MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0})) * $signed((taps_m_rsci_idat[351:341]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0 = $signed(delay_lane_m_0_sva)
      * $signed((taps_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0 = $signed(delay_lane_m_3_sva)
      * $signed((taps_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0 = $signed(delay_lane_m_4_sva)
      * $signed((taps_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0 = $signed(delay_lane_m_5_sva)
      * $signed((taps_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0 = $signed(delay_lane_m_6_sva)
      * $signed((taps_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0 = $signed(delay_lane_m_7_sva)
      * $signed((taps_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0 = $signed(delay_lane_m_8_sva)
      * $signed((taps_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0 = $signed(delay_lane_m_9_sva)
      * $signed((taps_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0 = $signed(delay_lane_m_10_sva)
      * $signed((taps_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0 = $signed(delay_lane_m_11_sva)
      * $signed((taps_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0 = $signed(delay_lane_m_12_sva)
      * $signed((taps_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0 = $signed(delay_lane_m_13_sva)
      * $signed((taps_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0 = $signed(delay_lane_m_14_sva)
      * $signed((taps_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0 = $signed(delay_lane_m_15_sva)
      * $signed((taps_m_rsci_idat[175:165]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0 = $signed(delay_lane_m_16_sva)
      * $signed((taps_m_rsci_idat[186:176]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0 = $signed(delay_lane_m_1_sva)
      * $signed((taps_m_rsci_idat[32:22]));
  assign nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = conv_s2s_5_6({MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4
      , MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0}) + 6'b000001;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:0];
  assign MAC_18_r_ac_float_else_and_nl = MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_18_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1
      = conv_s2s_6_7({MAC_18_r_ac_float_else_and_nl , MAC_18_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1[6:0];
  assign MAC_19_r_ac_float_else_and_nl = MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_19_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1
      = conv_s2s_6_7({MAC_19_r_ac_float_else_and_nl , MAC_19_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1[6:0];
  assign MAC_20_r_ac_float_else_and_nl = MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_20_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1
      = conv_s2s_6_7({MAC_20_r_ac_float_else_and_nl , MAC_20_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1[6:0];
  assign MAC_21_r_ac_float_else_and_nl = MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_21_r_ac_float_else_and_1_nl = MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      & MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_21_r_ac_float_else_and_2_nl = MUX_v_4_2_2(4'b0000, MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1,
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1
      = conv_s2s_6_7({MAC_21_r_ac_float_else_and_nl , MAC_21_r_ac_float_else_and_1_nl
      , MAC_21_r_ac_float_else_and_2_nl}) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1[6:0];
  assign MAC_22_r_ac_float_else_and_nl = MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_22_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1
      = conv_s2s_6_7({MAC_22_r_ac_float_else_and_nl , MAC_22_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1[6:0];
  assign MAC_23_r_ac_float_else_and_nl = MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_23_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1
      = conv_s2s_6_7({MAC_23_r_ac_float_else_and_nl , MAC_23_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1[6:0];
  assign MAC_24_r_ac_float_else_and_nl = MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_24_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1
      = conv_s2s_6_7({MAC_24_r_ac_float_else_and_nl , MAC_24_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1[6:0];
  assign MAC_25_r_ac_float_else_and_nl = MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_25_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1
      = conv_s2s_6_7({MAC_25_r_ac_float_else_and_nl , MAC_25_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1[6:0];
  assign MAC_26_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
      & MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_26_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0,
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1
      = conv_s2s_6_7({MAC_26_r_ac_float_else_and_nl , MAC_26_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1[6:0];
  assign MAC_27_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
      & MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_27_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0,
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1
      = conv_s2s_6_7({MAC_27_r_ac_float_else_and_nl , MAC_27_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1[6:0];
  assign MAC_28_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
      & MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_28_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0,
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1
      = conv_s2s_6_7({MAC_28_r_ac_float_else_and_nl , MAC_28_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1[6:0];
  assign MAC_29_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
      & MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_29_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0,
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1
      = conv_s2s_6_7({MAC_29_r_ac_float_else_and_nl , MAC_29_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1[6:0];
  assign MAC_30_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
      & MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_30_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0,
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1
      = conv_s2s_6_7({MAC_30_r_ac_float_else_and_nl , MAC_30_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1[6:0];
  assign MAC_31_r_ac_float_else_and_nl = MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_31_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1
      = conv_s2s_6_7({MAC_31_r_ac_float_else_and_nl , MAC_31_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1[6:0];
  assign MAC_1_r_ac_float_else_and_nl = MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_1_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1
      = conv_s2s_6_7({MAC_1_r_ac_float_else_and_nl , MAC_1_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[6:4])
      + 3'b001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign MAC_32_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
      & MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_32_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0,
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1 =
      conv_s2s_6_7({MAC_32_r_ac_float_else_and_nl , MAC_32_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1 = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[10]))
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[10])
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[10]))
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[10])
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[10]))
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[10])
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[10]))
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[10])
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[10]))
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[10])
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[10]))
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[10])
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0[10]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0[10])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0[10]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0[10])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0[10]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0[10])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0[10]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0[10])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0[10]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0[10])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10]))
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10])
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0[10]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0[10])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      =  -operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2)}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg)
      + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg)
      + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg)
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg)
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg)
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg)
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg)
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg)
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]))})
      + conv_u2s_5_7(MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)
      + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[4])})
      + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg)
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg)
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg)
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg)
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg)
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg)
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg)
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0[10]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0[10])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_18_sva_1[3:0];
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg) + 7'b0000001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0[10]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0[10])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_19_sva_1[3:0];
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg) + 7'b0000001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0[10]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0[10])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_20_sva_1[3:0];
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg) + 7'b0000001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0[10]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0[10])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_21_sva_1[3:0];
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg) + 7'b0000001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0[10]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0[10])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_22_sva_1[3:0];
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg) + 7'b0000001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0[10]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0[10])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_23_sva_1[3:0];
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg) + 7'b0000001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0[10]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0[10])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_24_sva_1[3:0];
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg) + 7'b0000001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0[10]))
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0[10])
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_25_sva_1[3:0];
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg) + 7'b0000001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[10]))
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[10])
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_26_sva_1[3:0];
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg) + 7'b0000001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[10]))
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[10])
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_27_sva_1[3:0];
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg) + 7'b0000001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[10]))
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[10])
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_28_sva_1[3:0];
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg) + 7'b0000001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[10]))
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[10])
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_29_sva_1[3:0];
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg) + 7'b0000001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[10]))
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[10])
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_30_sva_1[3:0];
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg) + 7'b0000001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[10]))
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[10])
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_31_sva_1[3:0];
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg) + 7'b0000001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[10]))
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[10])
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1[3:0];
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg) + 7'b0000001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3 = ~((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[5:4]==2'b01));
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      =  -(MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]);
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1])
      | nor_187_cse);
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6
      | nor_190_cse);
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6
      | nor_193_cse);
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6
      | nor_196_cse);
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6
      | nor_199_cse);
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
      | nor_202_cse);
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6
      | nor_207_cse);
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6
      | nor_210_cse);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6
      | nor_212_cse);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
      | nor_179_cse);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6
      | nor_177_cse);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6
      | nor_175_cse);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6
      | nor_173_cse);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6
      | nor_166_cse);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6
      | nor_164_cse);
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp
      = MUX1HOT_v_7_3_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp
      = MUX1HOT_v_7_3_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp
      = MUX1HOT_v_7_3_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp
      = MUX1HOT_v_7_3_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp
      = MUX1HOT_v_7_3_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp
      = MUX1HOT_v_7_3_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp
      = MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp
      = MUX1HOT_v_7_3_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp
      = MUX1HOT_v_7_3_2(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 + conv_u2s_4_7(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp
      = MUX1HOT_v_7_3_2(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 + conv_u2s_4_7(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp
      = MUX1HOT_v_7_3_2(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0)
      , (~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1)})
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp
      = MUX1HOT_v_7_3_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp
      = MUX1HOT_v_7_3_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[5:4]!=2'b00))));
  assign or_482_ssc = nor_169_cse | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0;
  assign MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4 = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1[0])
      & or_482_ssc;
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl = ~ or_482_ssc;
  assign MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0 = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      4'b1111, ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_1_lpi_1_dfm_1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl});
  assign nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl = conv_s2s_5_6({(~
      MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4) , (~ MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0)})
      + 6'b000001;
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl = nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl[5:0];
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1 =
      readslicef_6_1_5(MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 | nor_169_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4
      = MUX_v_2_2_2(2'b00, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4!=2'b00))));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_96_mx0
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm,
      MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva + conv_s2s_6_7({1'b1
      , (~ MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp
      = MUX1HOT_v_7_3_2(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[5:4]!=2'b00))));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_99_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_99_nl);
  assign nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      + conv_s2s_5_6({(~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0)
      , (~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1)})
      + 6'b000001;
  assign MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_3_result_operator_result_operator_nor_tmp = ~((result_m_1_lpi_1_dfm_1_10_7!=4'b0000)
      | result_m_1_lpi_1_dfm_1_6 | (result_m_1_lpi_1_dfm_1_5_4!=2'b00) | (result_m_1_lpi_1_dfm_1_3_0!=4'b0000));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7[3]) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7[3])
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign result_m_1_lpi_1_dfm_1_10_7 = MUX1HOT_v_4_3_2(4'b0111, 4'b1000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7,
      {result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp});
  assign result_m_1_lpi_1_dfm_1_6 = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc)) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_132_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_158_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_132_nl);
  assign result_m_1_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_158_nl,
      2'b11, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_133_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_159_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_133_nl);
  assign result_m_1_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_159_nl,
      4'b1111, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_32_ssc);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0);
  assign MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0);
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0);
  assign MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0);
  assign MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0);
  assign MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0);
  assign MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0);
  assign MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0);
  assign MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0);
  assign MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0);
  assign MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0);
  assign MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0);
  assign MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0);
  assign MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0);
  assign MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0);
  assign nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl
      = ({1'b1 , (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm)
      + 7'b0000001;
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl
      = nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl[6:0];
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1
      = readslicef_7_1_6(MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl);
  assign nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_s2s_5_6({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm)})
      + 6'b000001;
  assign MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[5:0];
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp
      = MUX_v_6_2_2(6'b110000, MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign or_tmp_1 = (~ (fsm_output[0])) | (fsm_output[7]);
  assign or_tmp_2 = (fsm_output[0]) | (fsm_output[7]);
  assign and_dcpl_1 = ~((fsm_output[7:6]!=2'b00));
  assign and_861_cse = (fsm_output[3:1]==3'b111);
  assign or_tmp_17 = (fsm_output[4]) | and_861_cse;
  assign nor_tmp_9 = (fsm_output[4:1]==4'b1111);
  assign or_tmp_25 = (fsm_output[1]) | (fsm_output[3]);
  assign and_tmp_3 = (fsm_output[6]) & or_tmp_25;
  assign nor_tmp_12 = (fsm_output[3]) & (fsm_output[6]);
  assign mux_tmp_73 = MUX_s_1_2_2((~ (fsm_output[0])), (fsm_output[0]), fsm_output[1]);
  assign or_tmp_62 = (fsm_output[1:0]!=2'b01);
  assign or_tmp_87 = (fsm_output[1:0]!=2'b00);
  assign and_dcpl_36 = ~((fsm_output[5:4]!=2'b00));
  assign or_dcpl_50 = (fsm_output[6]) | (fsm_output[2]) | or_359_cse;
  assign or_dcpl_54 = or_tmp_2 | or_tmp_25 | or_dcpl_50;
  assign or_dcpl_56 = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[4])))
      | (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[5]);
  assign and_dcpl_47 = ~((fsm_output[2]) | (fsm_output[4]));
  assign and_dcpl_48 = and_dcpl_47 & (~ (fsm_output[5]));
  assign and_dcpl_49 = (fsm_output[7]) & (fsm_output[0]);
  assign and_dcpl_50 = and_dcpl_49 & (~ (fsm_output[1]));
  assign and_dcpl_59 = ~((fsm_output[6]) | (fsm_output[2]));
  assign and_dcpl_60 = and_dcpl_59 & and_dcpl_36;
  assign and_dcpl_61 = ~((fsm_output[1]) | (fsm_output[3]));
  assign and_dcpl_63 = nor_66_cse & and_dcpl_61;
  assign and_dcpl_64 = and_dcpl_63 & and_dcpl_60;
  assign and_dcpl_65 = (fsm_output[1]) & (~ (fsm_output[3]));
  assign and_dcpl_66 = nor_66_cse & and_dcpl_65;
  assign and_dcpl_67 = and_dcpl_66 & and_dcpl_60;
  assign mux_tmp_110 = MUX_s_1_2_2(and_867_cse, nor_tmp_12, fsm_output[2]);
  assign or_tmp_92 = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]) | (fsm_output[1]);
  assign mux_tmp_113 = MUX_s_1_2_2(nor_tmp_12, and_tmp_3, fsm_output[2]);
  assign mux_tmp_116 = MUX_s_1_2_2(and_tmp_3, (fsm_output[6]), fsm_output[2]);
  assign not_tmp_115 = ~((fsm_output[6]) | (fsm_output[3]) | (fsm_output[1]));
  assign mux_tmp_119 = MUX_s_1_2_2(not_tmp_115, and_867_cse, fsm_output[2]);
  assign or_tmp_96 = (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[7]);
  assign or_tmp_100 = (fsm_output[1:0]!=2'b10);
  assign nor_tmp_24 = (fsm_output[3]) & (fsm_output[1]);
  assign mux_128_nl = MUX_s_1_2_2(and_dcpl_61, nor_tmp_24, fsm_output[6]);
  assign mux_tmp_126 = MUX_s_1_2_2(mux_128_nl, nor_tmp_12, fsm_output[2]);
  assign or_dcpl_66 = or_tmp_25 | (fsm_output[2]);
  assign or_tmp_102 = (fsm_output[4:1]!=4'b0000);
  assign mux_tmp_128 = MUX_s_1_2_2((~ or_tmp_102), nor_tmp_9, fsm_output[5]);
  assign mux_tmp_129 = MUX_s_1_2_2(nor_tmp_24, (fsm_output[3]), fsm_output[2]);
  assign and_tmp_6 = (fsm_output[4]) & mux_tmp_129;
  assign mux_tmp_131 = MUX_s_1_2_2((fsm_output[3]), or_tmp_25, fsm_output[2]);
  assign and_tmp_7 = (fsm_output[4]) & mux_tmp_131;
  assign and_tmp_8 = (fsm_output[4]) & or_dcpl_66;
  assign or_tmp_104 = (fsm_output[4]) | mux_tmp_129;
  assign or_tmp_105 = (fsm_output[4]) | mux_tmp_131;
  assign mux_tmp_136 = MUX_s_1_2_2((~ or_tmp_102), or_tmp_105, fsm_output[5]);
  assign mux_140_nl = MUX_s_1_2_2(and_dcpl_61, (fsm_output[3]), fsm_output[6]);
  assign mux_tmp_138 = MUX_s_1_2_2(mux_140_nl, and_tmp_3, fsm_output[2]);
  assign or_dcpl_68 = (~ (fsm_output[1])) | (fsm_output[3]);
  assign or_dcpl_71 = (~ (fsm_output[7])) | (fsm_output[0]) | or_dcpl_68 | or_dcpl_50;
  assign and_dcpl_89 = (~ (fsm_output[6])) & (fsm_output[2]);
  assign and_dcpl_90 = and_dcpl_89 & and_dcpl_36;
  assign and_dcpl_91 = and_dcpl_63 & and_dcpl_90;
  assign and_dcpl_93 = (~ (fsm_output[7])) & (fsm_output[0]);
  assign and_dcpl_95 = and_dcpl_93 & and_dcpl_65 & and_dcpl_60;
  assign and_dcpl_96 = ~((fsm_output[1:0]!=2'b00));
  assign or_dcpl_74 = or_165_cse | (fsm_output[2]);
  assign or_dcpl_75 = or_dcpl_74 | or_359_cse;
  assign and_dcpl_98 = and_dcpl_93 & (fsm_output[1]);
  assign and_dcpl_99 = or_dcpl_75 & and_dcpl_98;
  assign and_dcpl_100 = and_dcpl_93 & and_dcpl_61;
  assign and_dcpl_101 = and_dcpl_100 & and_dcpl_60;
  assign xor_dcpl_3 = (fsm_output[0]) ^ (fsm_output[1]);
  assign and_dcpl_103 = or_dcpl_75 & xor_dcpl_3 & (~ (fsm_output[7]));
  assign and_dcpl_104 = ~((fsm_output[7]) | (fsm_output[3]));
  assign nor_tmp_27 = (fsm_output[2]) & (fsm_output[6]) & (fsm_output[3]) & (fsm_output[1]);
  assign or_tmp_110 = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]) | and_880_cse;
  assign or_189_nl = (fsm_output[4]) | (fsm_output[2]);
  assign mux_tmp_145 = MUX_s_1_2_2(and_tmp_3, (fsm_output[6]), or_189_nl);
  assign not_tmp_131 = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3])
      | and_880_cse);
  assign mux_tmp_147 = MUX_s_1_2_2(mux_tmp_113, (fsm_output[6]), fsm_output[4]);
  assign mux_tmp_149 = MUX_s_1_2_2(mux_tmp_110, (fsm_output[6]), fsm_output[4]);
  assign mux_tmp_151 = MUX_s_1_2_2(nor_tmp_27, (fsm_output[6]), fsm_output[4]);
  assign and_tmp_9 = (fsm_output[4]) & mux_tmp_116;
  assign and_tmp_10 = (fsm_output[4]) & mux_tmp_113;
  assign and_tmp_11 = (fsm_output[4]) & mux_tmp_110;
  assign or_tmp_114 = (fsm_output[3]) | and_880_cse;
  assign and_dcpl_118 = and_dcpl_1 & (~ (fsm_output[5]));
  assign or_tmp_116 = (fsm_output[3:2]!=2'b00) | and_880_cse;
  assign or_dcpl_83 = or_tmp_1 | or_tmp_25 | or_dcpl_50;
  assign nor_tmp_29 = (fsm_output[4]) & (fsm_output[2]) & (fsm_output[6]) & (fsm_output[3])
      & (fsm_output[1]);
  assign and_dcpl_129 = xor_dcpl_3 & and_dcpl_104 & and_dcpl_60;
  assign and_dcpl_132 = (fsm_output[7]) & (~ (fsm_output[0])) & and_dcpl_65 & and_dcpl_60;
  assign and_dcpl_135 = nor_66_cse & (fsm_output[1]);
  assign and_dcpl_136 = and_dcpl_135 & nor_61_cse;
  assign and_dcpl_143 = and_dcpl_98 & nor_61_cse;
  assign and_dcpl_148 = and_dcpl_100 & and_dcpl_90;
  assign or_dcpl_89 = or_165_cse | or_359_cse;
  assign or_dcpl_96 = or_tmp_2 | or_dcpl_68 | or_dcpl_50;
  assign mux_169_nl = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_165_cse);
  assign or_219_nl = nor_61_cse | (fsm_output[7]);
  assign mux_170_nl = MUX_s_1_2_2(mux_169_nl, or_219_nl, fsm_output[2]);
  assign mux_171_nl = MUX_s_1_2_2(mux_170_nl, (fsm_output[7]), or_359_cse);
  assign and_dcpl_167 = (~ mux_171_nl) & and_dcpl_96;
  assign or_dcpl_100 = (fsm_output[7:6]!=2'b00);
  assign or_tmp_128 = (fsm_output[3]) | (~ or_tmp_100);
  assign and_dcpl_290 = and_dcpl_65 & (~ (fsm_output[6])) & and_dcpl_48;
  assign mux_203_nl = MUX_s_1_2_2(and_dcpl_61, or_tmp_25, fsm_output[6]);
  assign mux_tmp_201 = MUX_s_1_2_2(mux_203_nl, (fsm_output[6]), fsm_output[2]);
  assign and_dcpl_323 = nor_61_cse & (~ (fsm_output[2]));
  assign and_dcpl_324 = and_dcpl_323 & and_dcpl_36;
  assign and_dcpl_341 = (fsm_output[2]) & (~ (fsm_output[4]));
  assign and_dcpl_343 = not_tmp_115 & and_dcpl_341 & (~ (fsm_output[5]));
  assign and_dcpl_347 = nor_61_cse & (fsm_output[2]);
  assign and_dcpl_354 = (fsm_output[3]) & (~ (fsm_output[6]));
  assign and_dcpl_355 = and_dcpl_354 & (~ (fsm_output[2]));
  assign and_dcpl_360 = and_dcpl_354 & (fsm_output[2]);
  assign and_dcpl_365 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_382 = (fsm_output[5:4]==2'b10);
  assign and_dcpl_399 = (fsm_output[5:4]==2'b11);
  assign and_dcpl_416 = (~ (fsm_output[3])) & (fsm_output[6]);
  assign and_dcpl_417 = and_dcpl_416 & (~ (fsm_output[2]));
  assign and_dcpl_422 = and_dcpl_416 & (fsm_output[2]);
  assign and_dcpl_427 = nor_tmp_12 & (~ (fsm_output[2]));
  assign and_dcpl_432 = nor_tmp_12 & (fsm_output[2]);
  assign or_tmp_204 = (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]) | (~ or_tmp_100);
  assign or_dcpl_170 = or_dcpl_100 | or_359_cse;
  assign mux_tmp_284 = MUX_s_1_2_2((~ (fsm_output[1])), (fsm_output[1]), fsm_output[3]);
  assign mux_tmp_285 = MUX_s_1_2_2(mux_tmp_284, (fsm_output[3]), fsm_output[2]);
  assign and_dcpl_505 = and_dcpl_93 & (~ (fsm_output[1]));
  assign and_dcpl_514 = and_dcpl_59 & and_dcpl_365;
  assign and_dcpl_518 = and_dcpl_89 & and_dcpl_365;
  assign and_dcpl_524 = and_dcpl_135 & and_dcpl_354;
  assign and_dcpl_529 = and_dcpl_59 & and_dcpl_382;
  assign and_dcpl_533 = and_dcpl_89 & and_dcpl_382;
  assign and_dcpl_543 = and_dcpl_59 & and_dcpl_399;
  assign and_dcpl_547 = and_dcpl_89 & and_dcpl_399;
  assign and_dcpl_557 = (fsm_output[6]) & (~ (fsm_output[2]));
  assign and_dcpl_558 = and_dcpl_557 & and_dcpl_36;
  assign and_dcpl_564 = and_dcpl_135 & and_dcpl_416;
  assign and_dcpl_569 = (fsm_output[6]) & (fsm_output[2]);
  assign and_dcpl_570 = and_dcpl_569 & and_dcpl_36;
  assign and_dcpl_574 = and_dcpl_557 & and_dcpl_365;
  assign and_dcpl_578 = and_dcpl_569 & and_dcpl_365;
  assign and_dcpl_587 = and_dcpl_135 & nor_tmp_12;
  assign and_dcpl_589 = and_dcpl_557 & and_dcpl_382;
  assign and_dcpl_593 = and_dcpl_569 & and_dcpl_382;
  assign and_dcpl_609 = and_dcpl_557 & and_dcpl_399;
  assign and_dcpl_613 = and_dcpl_569 & and_dcpl_399;
  assign not_tmp_342 = ~((fsm_output[4]) | (fsm_output[2]) | (fsm_output[6]) | (fsm_output[3]));
  assign or_dcpl_180 = or_tmp_1 | or_dcpl_68 | or_dcpl_50;
  assign nor_tmp_33 = (fsm_output[6:5]==2'b11);
  assign or_495_cse = (fsm_output[4:3]!=2'b00);
  assign nor_tmp_36 = or_495_cse & (fsm_output[6:5]==2'b11);
  assign mux_tmp_351 = MUX_s_1_2_2(nor_203_cse, nor_tmp_33, or_495_cse);
  assign or_dcpl_200 = or_dcpl_100 | (fsm_output[5]);
  assign and_dcpl_688 = nor_66_cse & nor_tmp_24;
  assign and_dcpl_724 = and_dcpl_93 & (~ (fsm_output[1])) & (fsm_output[3]);
  assign return_e_rsci_idat_mx0c1 = and_dcpl_50 & nor_61_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & and_dcpl_48 & (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[5:4]==2'b01);
  assign operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 = or_tmp_87 &
      and_dcpl_104 & and_dcpl_60;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
      = and_dcpl_143 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
      = and_dcpl_143 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
      = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
      = and_dcpl_136 & and_dcpl_47 & (~((fsm_output[5]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3 = or_dcpl_89
      & and_dcpl_505;
  assign or_392_nl = (~ (fsm_output[3])) | (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_322_nl = MUX_s_1_2_2(or_392_nl, mux_420_cse, fsm_output[6]);
  assign mux_323_nl = MUX_s_1_2_2(mux_322_nl, mux_419_cse, fsm_output[2]);
  assign mux_324_nl = MUX_s_1_2_2(mux_323_nl, mux_416_cse, fsm_output[5]);
  assign mux_325_nl = MUX_s_1_2_2(mux_324_nl, mux_409_cse, fsm_output[4]);
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
      = (~ mux_325_nl) & and_dcpl_135;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
      = and_dcpl_135 & (fsm_output[3]) & (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_60;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
      = and_dcpl_135 & (fsm_output[3]) & (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_90;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_514;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_518;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7
      = and_dcpl_524 & (~ (fsm_output[2])) & (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_365;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
      = and_dcpl_135 & (fsm_output[3]) & (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_518;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_529;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_533;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
      = and_dcpl_135 & (fsm_output[3]) & (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_529;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
      = and_dcpl_135 & (fsm_output[3]) & (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_533;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_543;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_547;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
      = and_dcpl_135 & (fsm_output[3]) & (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_543;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
      = and_dcpl_135 & (fsm_output[3]) & (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_547;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_558;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
      = and_dcpl_564 & and_dcpl_341 & (~ (fsm_output[5])) & (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
      = and_dcpl_135 & (fsm_output[3]) & (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_558;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
      = and_dcpl_135 & (fsm_output[3]) & (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_570;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_574;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_578;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
      = and_dcpl_135 & (fsm_output[3]) & (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_574;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
      = and_dcpl_587 & (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[2]) & and_dcpl_365;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_589;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
      = and_dcpl_135 & (~ (fsm_output[3])) & (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_593;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
      = and_dcpl_587 & (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ (fsm_output[2])) & and_dcpl_382;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
      = and_dcpl_587 & (fsm_output[2]) & (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_382;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
      = and_dcpl_564 & (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ (fsm_output[2])) & and_dcpl_399;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
      = and_dcpl_564 & (fsm_output[2]) & (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_399;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
      = and_dcpl_135 & (fsm_output[3]) & (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_609;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32
      = and_dcpl_135 & (fsm_output[3]) & (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_613;
  assign or_tmp_270 = and_dcpl_688 | and_dcpl_66;
  assign and_tmp_15 = and_dcpl_66 & ((and_dcpl_514 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm)
      | (and_dcpl_518 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm)
      | (and_dcpl_529 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm)
      | (and_dcpl_547 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva)
      | (and_dcpl_533 & ac_float_cctor_operator_return_9_sva) | (and_dcpl_543 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva)
      | (and_dcpl_570 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva)
      | (and_dcpl_574 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva)
      | (and_dcpl_589 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm)
      | (and_dcpl_609 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
      & and_dcpl_613));
  assign or_tmp_283 = and_dcpl_688 | and_tmp_15;
  assign or_tmp_294 = (and_dcpl_514 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm)
      | (and_dcpl_518 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm)
      | (and_dcpl_529 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva)
      | (and_dcpl_547 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva)
      | (and_dcpl_533 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      | (and_dcpl_543 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva)
      | (and_dcpl_570 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva)
      | (and_dcpl_574 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva)
      | (and_dcpl_589 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (and_dcpl_609 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm)
      | (ac_float_cctor_operator_return_sva & and_dcpl_613);
  assign and_929_cse = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & and_dcpl_60;
  assign or_528_nl = and_929_cse | and_dcpl_66 | or_tmp_294;
  assign mux_tmp_427 = MUX_s_1_2_2(and_dcpl_66, or_528_nl, and_dcpl_688);
  assign nor_tmp_73 = (ac_float_cctor_operator_return_sva | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm)
      & and_dcpl_613;
  assign or_540_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | nor_tmp_73;
  assign mux_tmp_434 = MUX_s_1_2_2(nor_tmp_73, or_540_nl, and_dcpl_609);
  assign or_541_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
      | mux_tmp_434;
  assign mux_tmp_435 = MUX_s_1_2_2(mux_tmp_434, or_541_nl, and_dcpl_589);
  assign or_542_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      | mux_tmp_435;
  assign mux_tmp_436 = MUX_s_1_2_2(mux_tmp_435, or_542_nl, and_dcpl_574);
  assign or_543_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      | mux_tmp_436;
  assign mux_tmp_437 = MUX_s_1_2_2(mux_tmp_436, or_543_nl, and_dcpl_570);
  assign or_544_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_437;
  assign mux_tmp_438 = MUX_s_1_2_2(mux_tmp_437, or_544_nl, and_dcpl_543);
  assign or_545_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | ac_float_cctor_operator_return_9_sva | mux_tmp_438;
  assign mux_tmp_439 = MUX_s_1_2_2(mux_tmp_438, or_545_nl, and_dcpl_533);
  assign or_546_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | mux_tmp_439;
  assign mux_tmp_440 = MUX_s_1_2_2(mux_tmp_439, or_546_nl, and_dcpl_547);
  assign or_547_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | mux_tmp_440;
  assign mux_tmp_441 = MUX_s_1_2_2(mux_tmp_440, or_547_nl, and_dcpl_529);
  assign or_548_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | mux_tmp_441;
  assign mux_tmp_442 = MUX_s_1_2_2(mux_tmp_441, or_548_nl, and_dcpl_518);
  assign or_549_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_442;
  assign mux_446_nl = MUX_s_1_2_2(mux_tmp_442, or_549_nl, and_dcpl_514);
  assign mux_447_nl = MUX_s_1_2_2(or_tmp_294, mux_446_nl, and_dcpl_66);
  assign or_550_nl = and_929_cse | mux_447_nl;
  assign mux_tmp_445 = MUX_s_1_2_2(and_tmp_15, or_550_nl, and_dcpl_688);
  assign mux_449_nl = MUX_s_1_2_2(mux_tmp_445, mux_tmp_427, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign mux_436_nl = MUX_s_1_2_2(or_tmp_283, or_tmp_270, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign mux_450_nl = MUX_s_1_2_2(mux_449_nl, mux_436_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm);
  assign mux_tmp_448 = MUX_s_1_2_2(mux_tmp_445, mux_450_nl, and_dcpl_90);
  assign mux_470_nl = MUX_s_1_2_2(mux_tmp_427, or_tmp_270, and_cse);
  assign mux_452_nl = MUX_s_1_2_2(mux_tmp_448, mux_470_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva);
  assign mux_509_nl = MUX_s_1_2_2(or_tmp_283, or_tmp_270, and_901_cse);
  assign mux_435_nl = MUX_s_1_2_2(mux_509_nl, or_tmp_270, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva);
  assign mux_453_nl = MUX_s_1_2_2(mux_452_nl, mux_435_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign mux_tmp_451 = MUX_s_1_2_2(mux_tmp_448, mux_453_nl, and_dcpl_558);
  assign mux_508_nl = MUX_s_1_2_2(mux_tmp_427, or_tmp_270, and_cse);
  assign mux_432_nl = MUX_s_1_2_2(mux_508_nl, or_tmp_270, and_899_cse);
  assign mux_455_nl = MUX_s_1_2_2(mux_tmp_451, mux_432_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva);
  assign mux_471_nl = MUX_s_1_2_2(or_tmp_283, or_tmp_270, and_901_cse);
  assign mux_427_nl = MUX_s_1_2_2(mux_471_nl, or_tmp_270, and_902_cse);
  assign mux_434_nl = MUX_s_1_2_2(mux_427_nl, or_tmp_270, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva);
  assign mux_456_nl = MUX_s_1_2_2(mux_455_nl, mux_434_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign mux_tmp_454 = MUX_s_1_2_2(mux_tmp_451, mux_456_nl, and_dcpl_578);
  assign nor_294_cse = ~((fsm_output[1]) | (fsm_output[4]));
  assign nor_299_cse = ~((fsm_output[5]) | (fsm_output[3]));
  assign and_1120_cse = (~ (fsm_output[6])) & (fsm_output[2]) & nor_299_cse & nor_66_cse
      & nor_294_cse;
  assign and_352_ssc = nor_66_cse & (~ (fsm_output[1])) & (~(nor_169_cse | (fsm_output[3])))
      & and_dcpl_89 & (~ operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0)
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp & (fsm_output[5:4]==2'b00);
  assign and_358_ssc = (nor_169_cse | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0
      | (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp)) & nor_66_cse
      & and_dcpl_343;
  assign nor_30_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign mux_229_nl = MUX_s_1_2_2(or_tmp_62, mux_tmp_73, nor_30_nl);
  assign mux_230_nl = MUX_s_1_2_2(mux_229_nl, mux_tmp_73, MAC_3_result_operator_result_operator_nor_tmp);
  assign and_362_ssc = (~(mux_230_nl | (fsm_output[7]))) & and_dcpl_347 & and_dcpl_36;
  assign nor_171_nl = ~((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[4])));
  assign mux_257_nl = MUX_s_1_2_2(nor_171_nl, (fsm_output[4]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign or_327_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_326_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_256_nl = MUX_s_1_2_2(or_327_nl, or_326_nl, fsm_output[4]);
  assign mux_258_nl = MUX_s_1_2_2(mux_257_nl, mux_256_nl, fsm_output[2]);
  assign or_325_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_324_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_254_nl = MUX_s_1_2_2(or_325_nl, or_324_nl, fsm_output[4]);
  assign or_323_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_322_nl = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm;
  assign mux_253_nl = MUX_s_1_2_2(or_323_nl, or_322_nl, fsm_output[4]);
  assign mux_255_nl = MUX_s_1_2_2(mux_254_nl, mux_253_nl, fsm_output[2]);
  assign mux_259_nl = MUX_s_1_2_2(mux_258_nl, mux_255_nl, fsm_output[3]);
  assign or_321_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_320_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_250_nl = MUX_s_1_2_2(or_321_nl, or_320_nl, fsm_output[4]);
  assign or_319_nl = ac_float_cctor_operator_return_9_sva | (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_318_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_249_nl = MUX_s_1_2_2(or_319_nl, or_318_nl, fsm_output[4]);
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, mux_249_nl, fsm_output[2]);
  assign or_317_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_316_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_247_nl = MUX_s_1_2_2(or_317_nl, or_316_nl, fsm_output[4]);
  assign or_315_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_314_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_246_nl = MUX_s_1_2_2(or_315_nl, or_314_nl, fsm_output[4]);
  assign mux_248_nl = MUX_s_1_2_2(mux_247_nl, mux_246_nl, fsm_output[2]);
  assign mux_252_nl = MUX_s_1_2_2(mux_251_nl, mux_248_nl, fsm_output[3]);
  assign mux_260_nl = MUX_s_1_2_2(mux_259_nl, mux_252_nl, fsm_output[5]);
  assign or_313_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_312_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      | (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_242_nl = MUX_s_1_2_2(or_313_nl, or_312_nl, fsm_output[4]);
  assign or_311_nl = (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  assign or_310_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_241_nl = MUX_s_1_2_2(or_311_nl, or_310_nl, fsm_output[4]);
  assign mux_243_nl = MUX_s_1_2_2(mux_242_nl, mux_241_nl, fsm_output[2]);
  assign or_309_nl = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  assign or_308_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_239_nl = MUX_s_1_2_2(or_309_nl, or_308_nl, fsm_output[4]);
  assign or_307_nl = (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva;
  assign or_306_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
      | (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_238_nl = MUX_s_1_2_2(or_307_nl, or_306_nl, fsm_output[4]);
  assign mux_240_nl = MUX_s_1_2_2(mux_239_nl, mux_238_nl, fsm_output[2]);
  assign mux_244_nl = MUX_s_1_2_2(mux_243_nl, mux_240_nl, fsm_output[3]);
  assign or_305_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
      | (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_304_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_235_nl = MUX_s_1_2_2(or_305_nl, or_304_nl, fsm_output[4]);
  assign or_303_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
      | (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_302_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
      | (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_234_nl = MUX_s_1_2_2(or_303_nl, or_302_nl, fsm_output[4]);
  assign mux_236_nl = MUX_s_1_2_2(mux_235_nl, mux_234_nl, fsm_output[2]);
  assign or_301_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_300_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
      | (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_232_nl = MUX_s_1_2_2(or_301_nl, or_300_nl, fsm_output[4]);
  assign or_299_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_298_nl = ac_float_cctor_operator_return_sva | (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_231_nl = MUX_s_1_2_2(or_299_nl, or_298_nl, fsm_output[4]);
  assign mux_233_nl = MUX_s_1_2_2(mux_232_nl, mux_231_nl, fsm_output[2]);
  assign mux_237_nl = MUX_s_1_2_2(mux_236_nl, mux_233_nl, fsm_output[3]);
  assign mux_245_nl = MUX_s_1_2_2(mux_244_nl, mux_237_nl, fsm_output[5]);
  assign mux_261_nl = MUX_s_1_2_2(mux_260_nl, mux_245_nl, fsm_output[6]);
  assign and_365_ssc = mux_261_nl & nor_66_cse & (fsm_output[1]) & (~ MAC_3_result_operator_result_operator_nor_tmp);
  assign and_371_ssc = (((MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_355
      & and_dcpl_36;
  assign and_376_ssc = (((MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_360
      & and_dcpl_36;
  assign and_381_ssc = (((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_323
      & and_dcpl_365;
  assign and_385_ssc = (((MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_347
      & and_dcpl_365;
  assign and_389_ssc = (((MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_355
      & and_dcpl_365;
  assign and_393_ssc = (((MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_360
      & and_dcpl_365;
  assign and_398_ssc = (((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_323
      & and_dcpl_382;
  assign and_402_ssc = (((MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_9_sva)) | MAC_3_result_operator_result_operator_nor_tmp)
      & and_dcpl_135 & and_dcpl_347 & and_dcpl_382;
  assign and_406_ssc = (((MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_355
      & and_dcpl_382;
  assign and_410_ssc = (((MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_360
      & and_dcpl_382;
  assign and_415_ssc = (((MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_323
      & and_dcpl_399;
  assign and_419_ssc = (((MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_347
      & and_dcpl_399;
  assign and_423_ssc = (((MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_355
      & and_dcpl_399;
  assign and_427_ssc = (((MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_360
      & and_dcpl_399;
  assign and_433_ssc = (((MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_417
      & and_dcpl_36;
  assign and_438_ssc = (((MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_422
      & and_dcpl_36;
  assign and_443_ssc = (((MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_427
      & and_dcpl_36;
  assign and_448_ssc = (((MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_432
      & and_dcpl_36;
  assign and_452_ssc = (((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_417
      & and_dcpl_365;
  assign and_456_ssc = (((MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_422
      & and_dcpl_365;
  assign and_460_ssc = (((MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_427
      & and_dcpl_365;
  assign and_464_ssc = (((MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_432
      & and_dcpl_365;
  assign and_468_ssc = (((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_417
      & and_dcpl_382;
  assign and_472_ssc = (((MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_422
      & and_dcpl_382;
  assign and_476_ssc = (((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_427
      & and_dcpl_382;
  assign and_480_ssc = (((MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_432
      & and_dcpl_382;
  assign and_484_ssc = (((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_417
      & and_dcpl_399;
  assign and_488_ssc = (((MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_422
      & and_dcpl_399;
  assign and_492_ssc = (((MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_135 & and_dcpl_427
      & and_dcpl_399;
  assign and_496_ssc = (((MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_sva)) | MAC_3_result_operator_result_operator_nor_tmp)
      & and_dcpl_135 & and_dcpl_432 & and_dcpl_399;
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt = conv_s2s_5_6(delay_lane_e_9_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_itm
      = ~(and_dcpl_67 | ((or_dcpl_75 ^ (fsm_output[7])) & and_dcpl_96));
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0 = conv_s2s_5_6(delay_lane_e_10_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[54:50]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[5:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2}) + conv_s2s_6_7({1'b1
      , (~ MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg)}) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2}) + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl
      = MUX_v_7_2_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign and_898_nl = and_dcpl_67 & (~ or_553_tmp);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])))
      & and_dcpl_95;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_128_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])
      & and_dcpl_95;
  assign operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0 = MUX1HOT_v_7_5_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl,
      z_out_15, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      7'b1110000, {and_dcpl_101 , and_898_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_128_nl , or_553_tmp});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0
      = conv_s2s_5_6(delay_lane_e_25_sva) + conv_s2s_5_6(taps_e_rsci_idat[129:125]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0
      = conv_s2s_5_6(delay_lane_e_26_sva) + conv_s2s_5_6(taps_e_rsci_idat[134:130]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0
      = conv_s2s_5_6(delay_lane_e_27_sva) + conv_s2s_5_6(taps_e_rsci_idat[139:135]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0
      = conv_s2s_5_6(delay_lane_e_28_sva) + conv_s2s_5_6(taps_e_rsci_idat[144:140]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0
      = conv_s2s_5_6(delay_lane_e_0_sva) + conv_s2s_5_6(taps_e_rsci_idat[9:5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0
      = conv_s2s_5_6(delay_lane_e_29_sva) + conv_s2s_5_6(taps_e_rsci_idat[149:145]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0
      = conv_s2s_5_6({MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      , MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1})
      + conv_s2s_5_6(taps_e_rsci_idat[159:155]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0
      = conv_s2s_5_6(delay_lane_e_1_sva) + conv_s2s_5_6(taps_e_rsci_idat[14:10]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0
      = conv_s2s_5_6(delay_lane_e_3_sva) + conv_s2s_5_6(taps_e_rsci_idat[19:15]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0
      = conv_s2s_5_6(delay_lane_e_4_sva) + conv_s2s_5_6(taps_e_rsci_idat[24:20]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0
      = conv_s2s_5_6(delay_lane_e_5_sva) + conv_s2s_5_6(taps_e_rsci_idat[29:25]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0
      = conv_s2s_5_6(delay_lane_e_6_sva) + conv_s2s_5_6(taps_e_rsci_idat[34:30]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0
      = conv_s2s_5_6(delay_lane_e_7_sva) + conv_s2s_5_6(taps_e_rsci_idat[39:35]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0
      = conv_s2s_5_6(delay_lane_e_8_sva) + conv_s2s_5_6(taps_e_rsci_idat[44:40]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0[5:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc = and_dcpl_67
      | and_dcpl_95 | and_dcpl_99;
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_e_rsci_idat <= 5'b00000;
    end
    else if ( (and_dcpl_50 & and_dcpl_48 & or_dcpl_56 & nor_61_cse) | return_e_rsci_idat_mx0c1
        ) begin
      return_e_rsci_idat <= MUX_v_5_2_2((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[4:0]),
          5'b01111, return_e_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_m_rsci_idat <= 11'b00000000000;
    end
    else if ( ~((~((fsm_output[7]) & (fsm_output[0]))) | or_tmp_25 | or_dcpl_50)
        ) begin
      return_m_rsci_idat <= MUX1HOT_v_11_3_2(11'b01111111111, 11'b10000000000, (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:2]),
          {result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_31_nl
          , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse
        ) begin
      MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl,
          and_dcpl_67);
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_67);
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_67);
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_67);
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_67);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_67);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl,
          and_dcpl_67);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_54 ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      reg_return_e_triosy_obj_ld_cse <= 1'b0;
      reg_taps_e_triosy_obj_ld_cse <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= 18'b000000000000000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva <=
          4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1
          <= 2'b00;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0 <=
          1'b0;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1 <=
          4'b0000;
    end
    else begin
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0!=22'b0000000000000000000000);
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0!=22'b0000000000000000000000);
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0!=22'b0000000000000000000000);
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0!=22'b0000000000000000000000);
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0!=22'b0000000000000000000000);
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0!=22'b0000000000000000000000);
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0!=22'b0000000000000000000000);
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0!=22'b0000000000000000000000);
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0!=22'b0000000000000000000000);
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0!=22'b0000000000000000000000);
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0!=22'b0000000000000000000000);
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0!=22'b0000000000000000000000);
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0!=22'b0000000000000000000000);
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0!=22'b0000000000000000000000);
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0!=22'b0000000000000000000000);
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl,
          and_dcpl_67);
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl,
          and_dcpl_67);
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl,
          and_dcpl_67);
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl,
          and_dcpl_67);
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl,
          and_dcpl_67);
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl,
          and_dcpl_67);
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl,
          and_dcpl_67);
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
      reg_return_e_triosy_obj_ld_cse <= and_dcpl_49 & and_dcpl_61 & and_dcpl_60;
      reg_taps_e_triosy_obj_ld_cse <= ~ or_dcpl_54;
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[21:4];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_20_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_24_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_28_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= MUX_v_2_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl,
          and_dcpl_67);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm
          <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[3:0]),
          (z_out_16[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]),
          (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
          {and_163_nl , and_166_nl , and_169_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1
          <= MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm
          <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[3:0]),
          MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_14, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_15,
          {and_172_nl , and_175_nl , and_178_nl , and_dcpl_91 , and_dcpl_167});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1
          <= MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1
          <= MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1
          <= MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg[3:0]),
          MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_122_nl , and_185_nl , (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1
          <= MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg[3:0]),
          MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_123_nl , and_187_nl , (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva <=
          MUX1HOT_v_4_4_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[3:0]), (z_out_15[3:0]), {and_190_nl
          , and_193_nl , and_196_nl , and_dcpl_91});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg[3:0]),
          MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_125_nl , and_198_nl , (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[3:0]),
          MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_126_nl , and_200_nl , (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg[3:0]),
          MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_127_nl , and_202_nl , (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[3:0]),
          MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_128_nl , and_204_nl , (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[3:0]),
          MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_129_nl , and_206_nl , (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1
          <= MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[3:0]),
          MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_130_nl , and_208_nl , (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1
          <= MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg[3:0]),
          MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_131_nl , and_210_nl , (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1
          <= MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0 <=
          MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl,
          (MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4]), mux_127_itm);
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1 <=
          MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl,
          (MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[3:0]),
          mux_127_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_385_rgt | and_517_rgt ) begin
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[4:0]),
          {(~ and_76_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl
          , and_517_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_379_rgt | and_512_rgt ) begin
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0,
          {(~ nor_99_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl
          , and_512_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_372_rgt | and_507_rgt ) begin
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0,
          {(~ nor_100_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl
          , and_507_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_369_rgt | and_503_rgt ) begin
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0,
          {(~ nor_101_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl
          , and_503_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_363_rgt | and_499_rgt ) begin
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0,
          {(~ nor_102_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl
          , and_499_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_292_rgt | and_343_rgt ) begin
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0,
          {(~ nor_103_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl
          , and_343_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_281_rgt | and_333_rgt ) begin
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[4:0]),
          {(~ nor_104_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl
          , and_333_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_275_rgt | and_329_rgt ) begin
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[4:0]),
          {(~ and_85_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl
          , and_329_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_268_rgt | and_325_rgt ) begin
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[4:0]),
          {(~ and_87_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl
          , and_325_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_260_rgt | and_321_rgt ) begin
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[4:0]),
          {(~ and_89_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl
          , and_321_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_253_rgt | and_317_rgt ) begin
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[4:0]),
          {(~ and_91_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl
          , and_317_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_246_rgt | and_313_rgt ) begin
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[4:0]),
          {(~ and_92_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl
          , and_313_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_239_rgt | and_309_rgt ) begin
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[4:0]),
          {(~ and_93_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl
          , and_309_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_231_rgt | and_305_rgt ) begin
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[4:0]),
          {(~ and_94_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl
          , and_305_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_67 | or_287_rgt | and_339_rgt ) begin
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0,
          {(~ nor_105_rgt) , and_dcpl_67 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl
          , and_339_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_1_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_54 ) begin
      delay_lane_e_1_sva <= delay_lane_e_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_1_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      delay_lane_m_1_sva <= delay_lane_m_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_0_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_54 ) begin
      delay_lane_e_0_sva <= input_e_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_0_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_54 ) begin
      delay_lane_m_0_sva <= input_m_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_30_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_30_sva <= delay_lane_e_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_30_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_30_sva <= delay_lane_m_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_29_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_29_sva <= delay_lane_e_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_29_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_29_sva <= delay_lane_m_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_28_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_28_sva <= delay_lane_e_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_28_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_28_sva <= delay_lane_m_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_27_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_27_sva <= delay_lane_e_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_27_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_27_sva <= delay_lane_m_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_26_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_26_sva <= delay_lane_e_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_26_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_26_sva <= delay_lane_m_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_25_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_25_sva <= delay_lane_e_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_25_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_25_sva <= delay_lane_m_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_24_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_24_sva <= delay_lane_e_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_24_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_24_sva <= delay_lane_m_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_23_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_23_sva <= delay_lane_e_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_23_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_23_sva <= delay_lane_m_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_22_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_22_sva <= delay_lane_e_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_22_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_22_sva <= delay_lane_m_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_21_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_21_sva <= delay_lane_e_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_21_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_21_sva <= delay_lane_m_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_20_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_20_sva <= delay_lane_e_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_20_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_20_sva <= delay_lane_m_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_19_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_19_sva <= delay_lane_e_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_19_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_19_sva <= delay_lane_m_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_18_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_18_sva <= delay_lane_e_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_18_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_18_sva <= delay_lane_m_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_17_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_17_sva <= delay_lane_e_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_17_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_17_sva <= delay_lane_m_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_16_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_16_sva <= delay_lane_e_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_16_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_16_sva <= delay_lane_m_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_15_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_15_sva <= delay_lane_e_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_15_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_15_sva <= delay_lane_m_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_14_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_14_sva <= delay_lane_e_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_14_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_14_sva <= delay_lane_m_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_13_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_13_sva <= delay_lane_e_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_13_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_13_sva <= delay_lane_m_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_12_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_12_sva <= delay_lane_e_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_12_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_12_sva <= delay_lane_m_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_11_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_11_sva <= delay_lane_e_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_11_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_11_sva <= delay_lane_m_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_10_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_10_sva <= delay_lane_e_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_10_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_10_sva <= delay_lane_m_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_9_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_9_sva <= delay_lane_e_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_9_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_9_sva <= delay_lane_m_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_8_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_8_sva <= delay_lane_e_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_8_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_8_sva <= delay_lane_m_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_7_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_7_sva <= delay_lane_e_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_7_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_7_sva <= delay_lane_m_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_6_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_6_sva <= delay_lane_e_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_6_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_6_sva <= delay_lane_m_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_5_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_5_sva <= delay_lane_e_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_5_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_5_sva <= delay_lane_m_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_4_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_4_sva <= delay_lane_e_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_4_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_4_sva <= delay_lane_m_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_3_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_3_sva <= delay_lane_e_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_3_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_3_sva <= delay_lane_m_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_2_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_e_2_sva <= delay_lane_e_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_2_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_71 ) begin
      delay_lane_m_2_sva <= delay_lane_m_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
          <= 1'b0;
    end
    else if ( and_dcpl_64 | and_dcpl_67 | and_dcpl_91 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
          <= MUX1HOT_s_1_5_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[4]), (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
          (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
          {and_dcpl_64 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7 <= 4'b0000;
    end
    else if ( mux_505_nl & (~ (fsm_output[7])) ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7 <= MUX1HOT_v_4_49_2((z_out[12:9]),
          result_m_1_lpi_1_dfm_1_10_7, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_10_7,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10:7]),
          (z_out_1[12:9]), MAC_ac_float_cctor_m_4_lpi_1_dfm_10_7, (z_out_2[12:9]),
          MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7, (z_out_3[12:9]), MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7,
          (z_out_4[12:9]), MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7, (z_out_5[12:9]),
          MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7, (z_out_6[12:9]), MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7,
          (z_out_7[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[10:7]),
          (z_out_8[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[10:7]),
          (z_out_9[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[10:7]),
          (z_out_10[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[10:7]),
          (z_out_11[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[10:7]),
          (z_out_12[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[10:7]),
          (z_out_13[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[10:7]),
          (z_out_14[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[10:7]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10:7]),
          MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_26_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_27_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_28_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_29_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_30_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_31_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_lpi_1_dfm_10_7,
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[10:7]), {operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse , and_dcpl_99});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_371_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_209_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl
          , and_665_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_365_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_211_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_nl
          , and_661_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_361_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_213_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl
          , and_657_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_353_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_215_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_nl
          , and_653_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_347_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_217_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl
          , and_649_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_343_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_219_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_nl
          , and_645_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_339_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_221_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl
          , and_641_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_335_nl | (fsm_output[7]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_223_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0,
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_nl
          , and_637_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_390_nl & and_129_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_225_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_136_nl
          , and_689_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_387_nl & and_131_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_227_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl
          , and_685_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_384_nl & and_132_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_229_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl
          , and_681_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_381_nl & and_133_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_231_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_nl
          , and_677_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_378_nl & and_134_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_233_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_132_nl
          , and_673_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_374_nl) & and_135_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_235_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[4:0]),
          {and_dcpl_64 , and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl
          , and_669_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( and_dcpl_101 | and_dcpl_91 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= MUX_v_3_2_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp,
          and_dcpl_91);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_83 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva <= 7'b0000000;
    end
    else if ( ~(mux_165_nl & (~ (fsm_output[7])) & nor_61_cse & and_dcpl_36) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(((nor_187_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1]))
        & and_dcpl_98 & and_dcpl_324) | (~(mux_331_nl | (fsm_output[7])))) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_32_nl,
          5'b01111, {and_dcpl_101 , and_dcpl_67 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc ) begin
      MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7 <= MUX_v_4_2_2((z_out_17[10:7]), (delay_lane_m_30_sva[10:7]),
          and_dcpl_132);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc & (~ and_dcpl_67) ) begin
      MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0 <= MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (z_out_17[6:0]), (delay_lane_m_30_sva[6:0]), {and_dcpl_129 , and_dcpl_95
          , and_dcpl_132});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_26_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_27_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_28_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_29_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_30_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_31_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_4_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_lpi_1_dfm_10_7 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse ) begin
      MAC_ac_float_cctor_m_26_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_27_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_28_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_29_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_30_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_31_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_4_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1[10:7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse ) begin
      MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
      MAC_ac_float_cctor_m_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1[6:0]), and_dcpl_95);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
        | and_dcpl_148 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva <= MUX1HOT_v_11_5_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
          , and_dcpl_148});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= 1'b0;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
          <= MUX_s_1_2_2((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
          <= MUX_s_1_2_2((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
          <= MUX_s_1_2_2((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
          <= MUX_s_1_2_2((~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
          <= MUX_s_1_2_2((~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
          <= MUX_s_1_2_2((~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= MUX_s_1_2_2((~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= MUX_s_1_2_2((~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= MUX_s_1_2_2((~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= MUX_s_1_2_2((~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
          <= MUX_s_1_2_2((~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
          <= MUX_s_1_2_2((~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
          <= MUX_s_1_2_2((~ MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl,
          MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl,
          MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl,
          MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl,
          MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl,
          MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl,
          MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl,
          MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl,
          MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl,
          MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl,
          MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl,
          MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl,
          MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl,
          MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl,
          MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_95);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_96 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1
          <= MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= 1'b0;
    end
    else if ( and_dcpl_67 | and_dcpl_91 | and_dcpl_148 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= MUX1HOT_s_1_3_2((~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          (~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, {and_dcpl_67
          , and_dcpl_91 , and_dcpl_148});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= 1'b0;
    end
    else if ( and_dcpl_67 | and_dcpl_91 | and_dcpl_167 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= MUX1HOT_s_1_3_2((~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl,
          {and_dcpl_67 , and_dcpl_91 , and_dcpl_167});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva <= MUX1HOT_v_11_3_2((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva <= MUX1HOT_v_11_3_2((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva <= MUX1HOT_v_11_3_2((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva <= MUX1HOT_v_11_3_2((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva <= MUX1HOT_v_11_3_2((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva <= MUX1HOT_v_11_3_2((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva <= MUX1HOT_v_11_3_2((MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva <= MUX1HOT_v_11_3_2((MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva <= MUX1HOT_v_11_3_2((MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva <= MUX1HOT_v_11_3_2((MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva <= MUX1HOT_v_11_3_2((MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva <= MUX1HOT_v_11_3_2((MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva <= MUX1HOT_v_11_3_2((MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva <= MUX1HOT_v_11_3_2((MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
        | and_dcpl_95 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva <= MUX1HOT_v_11_3_2((MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
          , and_dcpl_95});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_96 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva[21]))
          & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp <= 1'b0;
    end
    else if ( and_dcpl_67 | and_dcpl_91 | and_dcpl_148 | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3
        ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_12, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl,
          result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3, {and_dcpl_67
          , and_dcpl_91 , and_dcpl_148 , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_10_7 <=
          4'b0000;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_6 <= 1'b0;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_5_4 <= 2'b00;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0 <= 4'b0000;
    end
    else if ( result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_10_7 <=
          MUX1HOT_v_4_32_2((z_out_17[10:7]), result_m_1_lpi_1_dfm_1_10_7, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10:7]),
          MAC_ac_float_cctor_m_4_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10:7]),
          MAC_ac_float_cctor_m_25_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_26_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_27_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_28_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_29_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_30_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_31_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_lpi_1_dfm_10_7,
          {and_dcpl_91 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_6 <= MUX1HOT_s_1_32_2((z_out_17[6]),
          result_m_1_lpi_1_dfm_1_6, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[6]),
          (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[6]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6]),
          {and_dcpl_91 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_5_4 <= MUX1HOT_v_2_32_2((z_out_17[5:4]),
          result_m_1_lpi_1_dfm_1_5_4, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[5:4]),
          (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[5:4]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[5:4]),
          {and_dcpl_91 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0 <= MUX1HOT_v_4_34_2((MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg[3:0]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (z_out_17[3:0]), result_m_1_lpi_1_dfm_1_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[3:0]),
          (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[3:0]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]),
          {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl , and_181_nl
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl , and_dcpl_91
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c32});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_180 ) begin
      ac_float_cctor_operator_return_sva <= ~((MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1!=11'b00000000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_9_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_180 ) begin
      ac_float_cctor_operator_return_9_sva <= ~((MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2!=11'b00000000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 2'b00;
    end
    else if ( and_dcpl_95 | and_dcpl_99 ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= MUX_v_2_2_2(MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          and_dcpl_99);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_67 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2
          <= 5'b00000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_itm
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
          <= MUX_s_1_2_2(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_32_nl,
          (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[5]),
          and_dcpl_101);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2
          <= MUX1HOT_v_5_5_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[4:0]),
          (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[4:0]),
          (z_out_16[4:0]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[4:0]),
          and_905_nl, {and_dcpl_64 , and_dcpl_95 , and_dcpl_99 , and_dcpl_101 , and_dcpl_103});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_or_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 <= MUX1HOT_s_1_50_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[6]),
          (z_out[8]), result_m_1_lpi_1_dfm_1_6, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_6,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[6]),
          (z_out_1[8]), (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[6]), (z_out_2[8]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6]), (z_out_3[8]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6]),
          (z_out_4[8]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6]), (z_out_5[8]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6]), (z_out_6[8]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6]),
          (z_out_7[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[6]),
          (z_out_8[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[6]),
          (z_out_9[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[6]),
          (z_out_10[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[6]),
          (z_out_11[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[6]),
          (z_out_12[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[6]),
          (z_out_13[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[6]),
          (z_out_14[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[6]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[6]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[6]), {operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1
          , operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse
          , and_dcpl_99});
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1 <= MUX1HOT_v_2_51_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[5:4]),
          (operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[5:4]), (z_out[7:6]),
          result_m_1_lpi_1_dfm_1_5_4, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_5_4,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[5:4]),
          (z_out_1[7:6]), (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[5:4]), (z_out_2[7:6]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[5:4]), (z_out_3[7:6]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[5:4]),
          (z_out_4[7:6]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[5:4]), (z_out_5[7:6]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[5:4]), (z_out_6[7:6]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[5:4]),
          (z_out_7[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[5:4]),
          (z_out_8[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[5:4]),
          (z_out_9[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[5:4]),
          (z_out_10[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[5:4]),
          (z_out_11[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[5:4]),
          (z_out_12[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[5:4]),
          (z_out_13[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[5:4]),
          (z_out_14[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[5:4]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[5:4]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[5:4]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[5:4]), {and_dcpl_64
          , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 , operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse , and_dcpl_99});
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 <= MUX1HOT_v_4_51_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[3:0]),
          (operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[3:0]), (z_out[5:2]),
          result_m_1_lpi_1_dfm_1_3_0, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_3_0,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[3:0]),
          (z_out_1[5:2]), (MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0[3:0]), (z_out_2[5:2]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]), (z_out_3[5:2]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]),
          (z_out_4[5:2]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]), (z_out_5[5:2]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]), (z_out_6[5:2]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]),
          (z_out_7[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_sva[3:0]),
          (z_out_8[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_sva[3:0]),
          (z_out_9[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_sva[3:0]),
          (z_out_10[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_sva[3:0]),
          (z_out_11[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_sva[3:0]),
          (z_out_12[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_sva[3:0]),
          (z_out_13[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_sva[3:0]),
          (z_out_14[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[3:0]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[3:0]),
          (MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[3:0]), {and_dcpl_64
          , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 , operator_13_2_true_AC_TRN_AC_WRAP_or_1_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_3_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_5_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_7_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_9_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_11_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_13_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse , operator_13_2_true_AC_TRN_AC_WRAP_or_15_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse , and_dcpl_99});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0 <= 8'b00000000;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 <= 4'b0000;
    end
    else if ( result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0 <= MUX_v_8_2_2((MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:4]),
          (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:4]),
          and_dcpl_99);
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl , and_183_nl
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl , and_dcpl_95
          , and_dcpl_99});
    end
  end
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_31_nl
      = ~((MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12]) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl = (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12])
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl
      = MUX_s_1_2_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl
      = MUX_s_1_2_2((MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg[4]), MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl
      = MUX_s_1_2_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl
      = MUX_s_1_2_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl
      = MUX_s_1_2_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_29_nl = MUX_s_1_2_2((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_29_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl = MUX_s_1_2_2((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_28_nl = MUX_s_1_2_2((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_28_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl = MUX_s_1_2_2((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_27_nl = MUX_s_1_2_2((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_27_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl = MUX_s_1_2_2((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_26_nl = MUX_s_1_2_2((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_20_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_26_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl = MUX_s_1_2_2((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_25_nl = MUX_s_1_2_2((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_25_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl = MUX_s_1_2_2((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_24_nl = MUX_s_1_2_2((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_24_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl = MUX_s_1_2_2((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_23_nl = MUX_s_1_2_2((MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_23_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl = MUX_s_1_2_2((MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_22_nl = MUX_s_1_2_2((MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_24_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_22_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl = MUX_s_1_2_2((MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_21_nl = MUX_s_1_2_2((MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_21_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl = MUX_s_1_2_2((MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_20_nl = MUX_s_1_2_2((MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_20_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl = MUX_s_1_2_2((MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_19_nl = MUX_s_1_2_2((MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_19_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl = MUX_s_1_2_2((MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_18_nl = MUX_s_1_2_2((MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_28_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_18_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl = MUX_s_1_2_2((MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_17_nl = MUX_s_1_2_2((MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_17_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl = MUX_s_1_2_2((MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_16_nl = MUX_s_1_2_2((MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_16_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_30_nl = MUX_s_1_2_2((MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_30_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_15_nl = MUX_v_2_2_2((MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:5]),
      (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl
      = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_15_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl
      = MUX_v_2_2_2(2'b00, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_seb);
  assign and_163_nl = and_dcpl_136 & and_dcpl_48 & (~((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_166_nl = and_dcpl_136 & and_dcpl_48 & (~ (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  assign and_169_nl = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign and_172_nl = and_dcpl_136 & and_dcpl_48 & (~((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_175_nl = and_dcpl_136 & and_dcpl_48 & (~ (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  assign and_178_nl = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]);
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_122_nl = ~(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_185_nl = MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_123_nl = ~(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_187_nl = MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign and_190_nl = and_dcpl_136 & and_dcpl_47 & (~ (fsm_output[5])) & (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]);
  assign and_193_nl = and_dcpl_136 & and_dcpl_48 & (~((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_196_nl = and_dcpl_136 & and_dcpl_48 & (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_25_lpi_1_dfm_6_0[3:0]);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_125_nl = ~(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_198_nl = MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_26_lpi_1_dfm_6_0[3:0]);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_126_nl = ~(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_200_nl = MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_27_lpi_1_dfm_6_0[3:0]);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_127_nl = ~(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_202_nl = MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_28_lpi_1_dfm_6_0[3:0]);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_128_nl = ~(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_204_nl = MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_29_lpi_1_dfm_6_0[3:0]);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_129_nl = ~(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_206_nl = MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_30_lpi_1_dfm_6_0[3:0]);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_130_nl = ~(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_208_nl = MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_31_lpi_1_dfm_6_0[3:0]);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_131_nl = ~(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_210_nl = MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_10_nl
      = MUX1HOT_s_1_35_2((MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4[0]),
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[4]),
      (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[4]),
      (MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4]),
      (delay_lane_e_30_sva[4]), {and_dcpl_67 , and_358_ssc , and_362_ssc , and_365_ssc
      , and_371_ssc , and_376_ssc , and_381_ssc , and_385_ssc , and_389_ssc , and_393_ssc
      , and_398_ssc , and_402_ssc , and_406_ssc , and_410_ssc , and_415_ssc , and_419_ssc
      , and_423_ssc , and_427_ssc , and_433_ssc , and_438_ssc , and_443_ssc , and_448_ssc
      , and_452_ssc , and_456_ssc , and_460_ssc , and_464_ssc , and_468_ssc , and_472_ssc
      , and_476_ssc , and_480_ssc , and_484_ssc , and_488_ssc , and_492_ssc , and_496_ssc
      , and_dcpl_132});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_10_nl
      & (~ and_352_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl
      = MUX_v_4_2_2(4'b0000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_16_nl
      = MUX1HOT_v_4_35_2((MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl,
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
      (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[3:0]),
      (MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]), (MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (delay_lane_e_30_sva[3:0]), {and_dcpl_67 , and_358_ssc , and_362_ssc , and_365_ssc
      , and_371_ssc , and_376_ssc , and_381_ssc , and_385_ssc , and_389_ssc , and_393_ssc
      , and_398_ssc , and_402_ssc , and_406_ssc , and_410_ssc , and_415_ssc , and_419_ssc
      , and_423_ssc , and_427_ssc , and_433_ssc , and_438_ssc , and_443_ssc , and_448_ssc
      , and_452_ssc , and_456_ssc , and_460_ssc , and_464_ssc , and_468_ssc , and_472_ssc
      , and_476_ssc , and_480_ssc , and_484_ssc , and_488_ssc , and_492_ssc , and_496_ssc
      , and_dcpl_132});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl
      = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_16_nl,
      4'b1111, and_352_ssc);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl = or_385_rgt & and_76_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl = or_379_rgt & nor_99_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl = or_372_rgt & nor_100_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl = or_369_rgt & nor_101_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl = or_363_rgt & nor_102_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl = or_292_rgt & nor_103_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl = or_281_rgt & nor_104_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl = or_275_rgt & and_85_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl = or_268_rgt & and_87_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl = or_260_rgt & and_89_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl = or_253_rgt & and_91_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl = or_246_rgt & and_92_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl = or_239_rgt & and_93_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl = or_231_rgt & and_94_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl = or_287_rgt & nor_105_rgt;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl = (~
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_67;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl =
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_67;
  assign or_568_nl = (~ (fsm_output[2])) | (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_499_nl = MUX_s_1_2_2((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_500_nl = MUX_s_1_2_2(or_568_nl, mux_499_nl, fsm_output[5]);
  assign mux_497_nl = MUX_s_1_2_2((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_496_nl = MUX_s_1_2_2((MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_498_nl = MUX_s_1_2_2(mux_497_nl, mux_496_nl, fsm_output[5]);
  assign mux_501_nl = MUX_s_1_2_2(mux_500_nl, mux_498_nl, fsm_output[4]);
  assign mux_493_nl = MUX_s_1_2_2((MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_492_nl = MUX_s_1_2_2((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_494_nl = MUX_s_1_2_2(mux_493_nl, mux_492_nl, fsm_output[5]);
  assign mux_490_nl = MUX_s_1_2_2((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_489_nl = MUX_s_1_2_2((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_491_nl = MUX_s_1_2_2(mux_490_nl, mux_489_nl, fsm_output[5]);
  assign mux_495_nl = MUX_s_1_2_2(mux_494_nl, mux_491_nl, fsm_output[4]);
  assign mux_502_nl = MUX_s_1_2_2(mux_501_nl, mux_495_nl, fsm_output[6]);
  assign mux_485_nl = MUX_s_1_2_2((MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_484_nl = MUX_s_1_2_2((MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_486_nl = MUX_s_1_2_2(mux_485_nl, mux_484_nl, fsm_output[5]);
  assign mux_482_nl = MUX_s_1_2_2((MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_481_nl = MUX_s_1_2_2((MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_483_nl = MUX_s_1_2_2(mux_482_nl, mux_481_nl, fsm_output[5]);
  assign mux_487_nl = MUX_s_1_2_2(mux_486_nl, mux_483_nl, fsm_output[4]);
  assign mux_478_nl = MUX_s_1_2_2((MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_477_nl = MUX_s_1_2_2((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, mux_477_nl, fsm_output[5]);
  assign mux_475_nl = MUX_s_1_2_2((MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_474_nl = MUX_s_1_2_2((MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]),
      (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]), fsm_output[2]);
  assign mux_476_nl = MUX_s_1_2_2(mux_475_nl, mux_474_nl, fsm_output[5]);
  assign mux_480_nl = MUX_s_1_2_2(mux_479_nl, mux_476_nl, fsm_output[4]);
  assign mux_488_nl = MUX_s_1_2_2(mux_487_nl, mux_480_nl, fsm_output[6]);
  assign mux_503_nl = MUX_s_1_2_2(mux_502_nl, mux_488_nl, fsm_output[3]);
  assign mux_504_nl = MUX_s_1_2_2(or_183_cse, (~ mux_503_nl), result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign and_1148_nl = (fsm_output[1]) & mux_504_nl;
  assign mux_505_nl = MUX_s_1_2_2(and_1148_nl, or_183_cse, fsm_output[0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl
      = ~((~ MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_nl
      = MUX1HOT_v_5_3_2((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_seb);
  assign or_437_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_4_0[4]);
  assign mux_366_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_437_nl);
  assign mux_367_nl = MUX_s_1_2_2(mux_366_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6);
  assign mux_368_nl = MUX_s_1_2_2((~ mux_367_nl), nor_tmp_27, fsm_output[4]);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, (fsm_output[6]), fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl = (mux_369_nl
      | (fsm_output[7])) & nor_106_ssc;
  assign and_665_nl = (nor_212_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_6)
      & and_dcpl_324 & nor_106_ssc;
  assign mux_370_nl = MUX_s_1_2_2(and_dcpl_323, nor_tmp_27, fsm_output[4]);
  assign mux_371_nl = MUX_s_1_2_2(mux_370_nl, (fsm_output[6]), fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      = ~((~ MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_nl
      = MUX1HOT_v_5_3_2((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_seb);
  assign or_433_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0[4]);
  assign mux_362_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_433_nl);
  assign mux_363_nl = MUX_s_1_2_2(mux_362_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6);
  assign nor_209_nl = ~((fsm_output[4]) | mux_363_nl);
  assign mux_364_nl = MUX_s_1_2_2(nor_209_nl, mux_tmp_145, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_nl = (mux_364_nl
      | (fsm_output[7])) & nor_107_ssc;
  assign and_661_nl = (nor_210_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_6)
      & and_dcpl_324 & nor_107_ssc;
  assign mux_365_nl = MUX_s_1_2_2(not_tmp_342, mux_tmp_145, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      = ~((~ MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_nl
      = MUX1HOT_v_5_3_2((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_seb);
  assign mux_359_nl = MUX_s_1_2_2(mux_tmp_351, nor_tmp_36, fsm_output[2]);
  assign or_428_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0[4]);
  assign mux_355_nl = MUX_s_1_2_2(nor_tmp_36, mux_tmp_351, or_428_nl);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, nor_tmp_36, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6);
  assign mux_357_nl = MUX_s_1_2_2(mux_tmp_351, mux_356_nl, fsm_output[0]);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, nor_tmp_33, fsm_output[2]);
  assign mux_360_nl = MUX_s_1_2_2(mux_359_nl, mux_358_nl, fsm_output[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl = (mux_360_nl
      | (fsm_output[7])) & nor_108_ssc;
  assign and_657_nl = (nor_207_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_6)
      & and_dcpl_324 & nor_108_ssc;
  assign mux_361_nl = MUX_s_1_2_2(not_tmp_342, mux_tmp_147, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      = ~((~ MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_nl
      = MUX1HOT_v_5_3_2((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_seb);
  assign nor_201_nl = ~((fsm_output[3]) | (fsm_output[5]) | (fsm_output[6]));
  assign nor_204_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6
      | nor_202_cse | (fsm_output[6:5]!=2'b00));
  assign mux_348_nl = MUX_s_1_2_2(nor_203_cse, nor_204_nl, fsm_output[0]);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, nor_tmp_33, fsm_output[3]);
  assign mux_350_nl = MUX_s_1_2_2(nor_201_nl, mux_349_nl, fsm_output[1]);
  assign and_882_nl = (fsm_output[3]) & (fsm_output[5]) & (fsm_output[6]);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, and_882_nl, fsm_output[2]);
  assign mux_352_nl = MUX_s_1_2_2(mux_351_nl, nor_tmp_33, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_nl = (mux_352_nl
      | (fsm_output[7])) & nor_109_ssc;
  assign and_653_nl = (nor_202_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_6)
      & and_dcpl_324 & nor_109_ssc;
  assign mux_353_nl = MUX_s_1_2_2(not_tmp_342, mux_tmp_149, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl
      = ~((~ MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_nl
      = MUX1HOT_v_5_3_2((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_seb);
  assign or_416_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0[4]);
  assign mux_344_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_416_nl);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6);
  assign nor_198_nl = ~((fsm_output[4]) | mux_345_nl);
  assign mux_346_nl = MUX_s_1_2_2(nor_198_nl, mux_tmp_151, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl = (mux_346_nl
      | (fsm_output[7])) & nor_110_ssc;
  assign and_649_nl = (nor_199_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_6)
      & and_dcpl_324 & nor_110_ssc;
  assign mux_347_nl = MUX_s_1_2_2(not_tmp_342, mux_tmp_151, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      = ~((~ MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_nl
      = MUX1HOT_v_5_3_2((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_seb);
  assign or_412_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0[4]);
  assign mux_340_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_412_nl);
  assign mux_341_nl = MUX_s_1_2_2(mux_340_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6);
  assign nor_195_nl = ~((fsm_output[4]) | mux_341_nl);
  assign mux_342_nl = MUX_s_1_2_2(nor_195_nl, and_tmp_9, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_nl = (mux_342_nl
      | (fsm_output[7])) & nor_111_ssc;
  assign and_645_nl = (nor_196_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_6)
      & and_dcpl_324 & nor_111_ssc;
  assign mux_343_nl = MUX_s_1_2_2(not_tmp_342, and_tmp_9, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl
      = ~((~ MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_nl
      = MUX1HOT_v_5_3_2((MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_seb);
  assign or_408_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0[4]);
  assign mux_336_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_408_nl);
  assign mux_337_nl = MUX_s_1_2_2(mux_336_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6);
  assign nor_192_nl = ~((fsm_output[4]) | mux_337_nl);
  assign mux_338_nl = MUX_s_1_2_2(nor_192_nl, and_tmp_10, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl = (mux_338_nl
      | (fsm_output[7])) & nor_112_ssc;
  assign and_641_nl = (nor_193_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_6)
      & and_dcpl_324 & nor_112_ssc;
  assign mux_339_nl = MUX_s_1_2_2(not_tmp_342, and_tmp_10, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      = ~((~ MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_nl
      = MUX1HOT_v_5_3_2((MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_seb);
  assign or_404_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0[4]);
  assign mux_332_nl = MUX_s_1_2_2(or_tmp_110, or_dcpl_74, or_404_nl);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, or_tmp_110, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6);
  assign nor_189_nl = ~((fsm_output[4]) | mux_333_nl);
  assign mux_334_nl = MUX_s_1_2_2(nor_189_nl, and_tmp_11, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_nl = (mux_334_nl
      | (fsm_output[7])) & nor_113_ssc;
  assign and_637_nl = (nor_190_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_6)
      & and_dcpl_324 & nor_113_ssc;
  assign mux_335_nl = MUX_s_1_2_2(not_tmp_342, and_tmp_11, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl
      = ~((~ MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_nl
      = MUX1HOT_v_5_3_2((MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_seb);
  assign or_478_nl = (fsm_output[3]) | ((nor_231_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[6]))
      & (fsm_output[1:0]==2'b11));
  assign mux_388_nl = MUX_s_1_2_2(or_tmp_114, or_478_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm);
  assign mux_389_nl = MUX_s_1_2_2((~ mux_388_nl), nor_tmp_24, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_136_nl = (mux_389_nl
      | or_dcpl_170) & and_129_ssc;
  assign and_689_nl = (nor_231_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm))
      & and_dcpl_290 & and_129_ssc;
  assign mux_390_nl = MUX_s_1_2_2((fsm_output[3]), (~ nor_tmp_24), fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl
      = ~((~ MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_nl
      = MUX1HOT_v_5_3_2((MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_seb);
  assign or_471_nl = (fsm_output[3]) | ((nor_227_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[6]))
      & (fsm_output[1:0]==2'b11));
  assign mux_385_nl = MUX_s_1_2_2(or_tmp_114, or_471_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign nor_229_nl = ~((fsm_output[2]) | mux_385_nl);
  assign mux_386_nl = MUX_s_1_2_2(nor_229_nl, or_dcpl_66, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl = (mux_386_nl
      | or_dcpl_200) & and_131_ssc;
  assign and_685_nl = (nor_227_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm))
      & and_dcpl_290 & and_131_ssc;
  assign mux_387_nl = MUX_s_1_2_2(or_92_cse, (~ or_dcpl_66), fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl
      = ~((~ MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_nl
      = MUX1HOT_v_5_3_2((MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_seb);
  assign or_464_nl = (fsm_output[3]) | ((nor_223_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[6]))
      & (fsm_output[1:0]==2'b11));
  assign mux_382_nl = MUX_s_1_2_2(or_tmp_114, or_464_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign nor_225_nl = ~((fsm_output[2]) | mux_382_nl);
  assign mux_383_nl = MUX_s_1_2_2(nor_225_nl, mux_tmp_131, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl = (mux_383_nl
      | or_dcpl_200) & and_132_ssc;
  assign and_681_nl = (nor_223_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm))
      & and_dcpl_290 & and_132_ssc;
  assign mux_384_nl = MUX_s_1_2_2(or_92_cse, (~ mux_tmp_131), fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl
      = ~((~ MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_nl
      = MUX1HOT_v_5_3_2((MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_seb);
  assign or_457_nl = (fsm_output[3]) | ((nor_219_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[6]))
      & (fsm_output[1:0]==2'b11));
  assign mux_379_nl = MUX_s_1_2_2(or_tmp_114, or_457_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign nor_221_nl = ~((fsm_output[2]) | mux_379_nl);
  assign mux_380_nl = MUX_s_1_2_2(nor_221_nl, mux_tmp_129, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_nl = (mux_380_nl
      | or_dcpl_200) & and_133_ssc;
  assign and_677_nl = (nor_219_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm))
      & and_dcpl_290 & and_133_ssc;
  assign mux_381_nl = MUX_s_1_2_2(or_92_cse, (~ mux_tmp_129), fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl
      = ~((~ MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_nl
      = MUX1HOT_v_5_3_2((MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_seb);
  assign or_450_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[5:4]!=2'b00);
  assign mux_375_nl = MUX_s_1_2_2(or_tmp_116, or_92_cse, or_450_nl);
  assign or_449_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[6]);
  assign mux_376_nl = MUX_s_1_2_2(mux_375_nl, or_tmp_116, or_449_nl);
  assign mux_377_nl = MUX_s_1_2_2((~ mux_376_nl), and_861_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_132_nl = (mux_377_nl
      | or_dcpl_200) & and_134_ssc;
  assign and_673_nl = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm))
      & and_dcpl_290 & and_134_ssc;
  assign mux_378_nl = MUX_s_1_2_2(or_92_cse, (~ and_861_cse), fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl
      = ~((~ MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_nl
      = MUX1HOT_v_5_3_2((MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_seb);
  assign or_443_nl = (fsm_output[3]) | ((nor_214_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6]))
      & (fsm_output[1:0]==2'b11));
  assign mux_372_nl = MUX_s_1_2_2(or_tmp_114, or_443_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign nor_216_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_372_nl);
  assign mux_373_nl = MUX_s_1_2_2(nor_216_nl, or_tmp_102, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl = (mux_373_nl
      | or_dcpl_100) & and_135_ssc;
  assign and_669_nl = (nor_214_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm))
      & and_dcpl_290 & and_135_ssc;
  assign nor_93_nl = ~((fsm_output[4:2]!=3'b000));
  assign mux_374_nl = MUX_s_1_2_2(nor_93_nl, or_tmp_102, fsm_output[5]);
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[2:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_18_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_19_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_20_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_21_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_22_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_23_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_24_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_25_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_26_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_27_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_28_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_29_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_30_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_31_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:4])
      + 3'b001;
  assign MAC_3_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_5
      & MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_3_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_4_0,
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva 
      = conv_s2s_6_7({MAC_3_r_ac_float_else_and_nl , MAC_3_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign mux_165_nl = MUX_s_1_2_2((fsm_output[1]), (~ or_tmp_87), fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl
      = ~((~ MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_nl
      = MUX1HOT_v_5_3_2((MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_32_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_seb);
  assign mux_166_nl = MUX_s_1_2_2(not_tmp_131, nor_tmp_29, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl
      = ~(mux_166_nl | (fsm_output[7]));
  assign mux_331_nl = MUX_s_1_2_2(not_tmp_342, nor_tmp_29, fsm_output[5]);
  assign MAC_11_r_ac_float_else_and_nl = MUX_v_2_2_2(2'b00, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1,
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign MAC_11_r_ac_float_else_and_1_nl = MUX_v_4_2_2(4'b0000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_11_r_ac_float_else_and_nl , MAC_11_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_12_r_ac_float_else_and_nl = MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_12_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_12_r_ac_float_else_and_nl , MAC_12_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_13_r_ac_float_else_and_nl = MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_13_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_13_r_ac_float_else_and_nl , MAC_13_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_14_r_ac_float_else_and_nl = MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_14_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_14_r_ac_float_else_and_nl , MAC_14_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_15_r_ac_float_else_and_nl = MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_15_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_15_r_ac_float_else_and_nl , MAC_15_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_16_r_ac_float_else_and_nl = MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_16_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_16_r_ac_float_else_and_nl , MAC_16_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_17_r_ac_float_else_and_nl = MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_17_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_17_r_ac_float_else_and_nl , MAC_17_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_2_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_5
      & MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_2_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_4_0,
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_2_r_ac_float_else_and_nl , MAC_2_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_4_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_5
      & MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_4_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_4_0,
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_4_r_ac_float_else_and_nl , MAC_4_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_5_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_5
      & MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_5_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_4_0,
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_5_r_ac_float_else_and_nl , MAC_5_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_6_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_5
      & MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_6_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_4_0,
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_6_r_ac_float_else_and_nl , MAC_6_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_7_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_5
      & MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_7_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_4_0,
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_7_r_ac_float_else_and_nl , MAC_7_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_8_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_5
      & MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_8_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_4_0,
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_8_r_ac_float_else_and_nl , MAC_8_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_9_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_5
      & MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_9_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_4_0,
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_9_r_ac_float_else_and_nl , MAC_9_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva[21]))
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva[21]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva[21]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva[21]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva[21]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva[21]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva[21]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva[21]))
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm);
  assign MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva[21]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva[21]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva[21]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva[21]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva[21]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva[21]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4!=11'b00000000000));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_13 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva[21]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl
      = ~((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1[5:4]==2'b01));
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl = ((~(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])))
      & and_dcpl_67) | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_11_itm_mx0c7;
  assign and_181_nl = MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & and_dcpl_67;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl = (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_67;
  assign nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:4])
      + 2'b01;
  assign MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (z_out_16[5:4]) + 2'b01;
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_32_nl = MUX1HOT_s_1_3_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[5]),
      (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5]), (z_out_16[5]),
      {and_dcpl_64 , and_dcpl_95 , and_dcpl_99});
  assign nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign and_696_nl = and_dcpl_505 & (fsm_output[5:3]==3'b000) & (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp
      | (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[5:4]!=2'b01))
      & and_dcpl_89;
  assign nand_18_nl = ~((fsm_output[1]) & or_183_cse);
  assign or_502_nl = (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp &
      (fsm_output[2])) | (fsm_output[6:3]!=4'b0000);
  assign nor_237_nl = ~((~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp)
      | (fsm_output[6:2]!=5'b00001));
  assign mux_391_nl = MUX_s_1_2_2(or_502_nl, nor_237_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign mux_392_nl = MUX_s_1_2_2(or_183_cse, mux_391_nl, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[4]);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, or_183_cse, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_128_tmp[5]);
  assign or_489_nl = (fsm_output[1]) | (~ mux_393_nl);
  assign mux_394_nl = MUX_s_1_2_2(nand_18_nl, or_489_nl, fsm_output[0]);
  assign or_555_nl = mux_394_nl | (fsm_output[7]);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_96_nl = (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_698_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_97_nl = (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_698_m1c & (~ mux_461_tmp);
  assign and_701_nl = or_dcpl_89 & (~ (fsm_output[7])) & or_dcpl_56 & (~ or_tmp_62);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_98_nl = (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_703_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_99_nl = (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_703_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_100_nl = (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_704_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_101_nl = (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_704_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_102_nl = (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_705_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_103_nl = (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_705_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_104_nl = (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_706_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_105_nl = (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_706_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_106_nl = (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_707_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_107_nl = (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_707_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_108_nl = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_708_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_109_nl = (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_708_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_110_nl = (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_709_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_111_nl = (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_709_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_112_nl = (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_710_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_113_nl = (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_710_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_114_nl = (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_711_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_115_nl = (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_711_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_116_nl = (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_712_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_117_nl = (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_712_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_118_nl = (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_713_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_119_nl = (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_713_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_120_nl = (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_714_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_121_nl = (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_714_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_122_nl = (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_715_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_123_nl = (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_715_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_124_nl = (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_716_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_125_nl = (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_716_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_126_nl = (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_717_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl = (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_717_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_nl = (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_718_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_129_nl = (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_718_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_130_nl = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_719_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_131_nl = (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_719_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_132_nl = (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_720_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_133_nl = (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_720_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_134_nl = (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_721_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_135_nl = (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_721_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_136_nl = (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_722_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_137_nl = (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_722_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_138_nl = (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_723_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_139_nl = (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_723_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_140_nl = (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_724_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_141_nl = (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_724_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_142_nl = (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_725_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_143_nl = (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_725_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_144_nl = (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_726_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_145_nl = (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_726_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_146_nl = (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_727_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_147_nl = (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_727_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_148_nl = (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_728_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_149_nl = (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_728_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_150_nl = (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_729_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_151_nl = (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_729_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_152_nl = (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_730_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_153_nl = (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_730_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_154_nl = (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_731_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_155_nl = (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_731_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_156_nl = (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_732_m1c & (~ mux_461_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_157_nl = (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_732_m1c & (~ mux_461_tmp);
  assign mux1h_1_nl = MUX1HOT_v_5_65_2((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1[4:0]),
      5'b01111, (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[4:0]),
      (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, {and_696_nl
      , or_555_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_96_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_97_nl
      , and_701_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_98_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_99_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_100_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_101_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_102_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_103_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_104_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_105_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_106_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_107_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_108_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_109_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_110_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_111_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_112_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_113_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_114_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_115_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_116_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_117_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_118_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_119_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_120_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_121_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_122_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_123_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_124_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_125_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_126_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_129_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_130_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_131_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_132_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_133_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_134_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_135_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_136_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_137_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_138_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_139_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_140_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_141_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_142_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_143_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_144_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_145_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_146_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_147_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_148_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_149_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_150_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_151_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_152_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_153_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_154_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_155_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_156_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_157_nl});
  assign not_995_nl = ~ mux_461_tmp;
  assign and_905_nl = MUX_v_5_2_2(5'b00000, mux1h_1_nl, not_995_nl);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl = (~(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])))
      & and_dcpl_67;
  assign and_183_nl = MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & and_dcpl_67;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl = (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_67;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl
      = MUX_v_7_2_2(MAC_ac_float_cctor_m_4_lpi_1_dfm_6_0, (signext_7_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]))),
      and_1120_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl
      = ~(and_1120_cse & (~(and_dcpl_59 & nor_299_cse & (~ (fsm_output[7])) & (fsm_output[0])
      & (fsm_output[1]) & (~ (fsm_output[4])))));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      = MUX_v_5_2_2((~ MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0),
      5'b00001, and_1120_cse);
  assign nl_acc_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl})
      + conv_s2u_7_8({(~ and_1120_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[7:0];
  assign z_out_15 = readslicef_8_7_1(acc_nl);
  assign and_1151_nl = or_183_cse & (~ (fsm_output[7])) & (fsm_output[0]) & (fsm_output[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl
      = MUX_v_5_2_2((signext_5_4(~ (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]))),
      ({MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      , MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1}),
      and_1151_nl);
  assign nl_z_out_16 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl)
      + 6'b000001;
  assign z_out_16 = nl_z_out_16[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_m1c = MUX_s_1_2_2((~
      MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1),
      (~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1),
      and_1120_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl = (~ and_1120_cse)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_m1c;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl = and_1120_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_m1c;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_158_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[10]))
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_159_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_158_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_159_nl, and_1120_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_160_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva[10])
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_160_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_nl, and_1120_cse);
  assign z_out_17 = MUX1HOT_v_11_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_sva,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva, 11'b01111111111,
      11'b10000000000, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl});

  function automatic  MUX1HOT_s_1_32_2;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [31:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    MUX1HOT_s_1_32_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_35_2;
    input  input_34;
    input  input_33;
    input  input_32;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [34:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    result = result | (input_32 & sel[32]);
    result = result | (input_33 & sel[33]);
    result = result | (input_34 & sel[34]);
    MUX1HOT_s_1_35_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_50_2;
    input  input_49;
    input  input_48;
    input  input_47;
    input  input_46;
    input  input_45;
    input  input_44;
    input  input_43;
    input  input_42;
    input  input_41;
    input  input_40;
    input  input_39;
    input  input_38;
    input  input_37;
    input  input_36;
    input  input_35;
    input  input_34;
    input  input_33;
    input  input_32;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [49:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    result = result | (input_32 & sel[32]);
    result = result | (input_33 & sel[33]);
    result = result | (input_34 & sel[34]);
    result = result | (input_35 & sel[35]);
    result = result | (input_36 & sel[36]);
    result = result | (input_37 & sel[37]);
    result = result | (input_38 & sel[38]);
    result = result | (input_39 & sel[39]);
    result = result | (input_40 & sel[40]);
    result = result | (input_41 & sel[41]);
    result = result | (input_42 & sel[42]);
    result = result | (input_43 & sel[43]);
    result = result | (input_44 & sel[44]);
    result = result | (input_45 & sel[45]);
    result = result | (input_46 & sel[46]);
    result = result | (input_47 & sel[47]);
    result = result | (input_48 & sel[48]);
    result = result | (input_49 & sel[49]);
    MUX1HOT_s_1_50_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_4_2;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [3:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    MUX1HOT_v_11_4_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_5_2;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [4:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    MUX1HOT_v_11_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_32_2;
    input [1:0] input_31;
    input [1:0] input_30;
    input [1:0] input_29;
    input [1:0] input_28;
    input [1:0] input_27;
    input [1:0] input_26;
    input [1:0] input_25;
    input [1:0] input_24;
    input [1:0] input_23;
    input [1:0] input_22;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [31:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    result = result | (input_22 & {2{sel[22]}});
    result = result | (input_23 & {2{sel[23]}});
    result = result | (input_24 & {2{sel[24]}});
    result = result | (input_25 & {2{sel[25]}});
    result = result | (input_26 & {2{sel[26]}});
    result = result | (input_27 & {2{sel[27]}});
    result = result | (input_28 & {2{sel[28]}});
    result = result | (input_29 & {2{sel[29]}});
    result = result | (input_30 & {2{sel[30]}});
    result = result | (input_31 & {2{sel[31]}});
    MUX1HOT_v_2_32_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_51_2;
    input [1:0] input_50;
    input [1:0] input_49;
    input [1:0] input_48;
    input [1:0] input_47;
    input [1:0] input_46;
    input [1:0] input_45;
    input [1:0] input_44;
    input [1:0] input_43;
    input [1:0] input_42;
    input [1:0] input_41;
    input [1:0] input_40;
    input [1:0] input_39;
    input [1:0] input_38;
    input [1:0] input_37;
    input [1:0] input_36;
    input [1:0] input_35;
    input [1:0] input_34;
    input [1:0] input_33;
    input [1:0] input_32;
    input [1:0] input_31;
    input [1:0] input_30;
    input [1:0] input_29;
    input [1:0] input_28;
    input [1:0] input_27;
    input [1:0] input_26;
    input [1:0] input_25;
    input [1:0] input_24;
    input [1:0] input_23;
    input [1:0] input_22;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [50:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    result = result | (input_22 & {2{sel[22]}});
    result = result | (input_23 & {2{sel[23]}});
    result = result | (input_24 & {2{sel[24]}});
    result = result | (input_25 & {2{sel[25]}});
    result = result | (input_26 & {2{sel[26]}});
    result = result | (input_27 & {2{sel[27]}});
    result = result | (input_28 & {2{sel[28]}});
    result = result | (input_29 & {2{sel[29]}});
    result = result | (input_30 & {2{sel[30]}});
    result = result | (input_31 & {2{sel[31]}});
    result = result | (input_32 & {2{sel[32]}});
    result = result | (input_33 & {2{sel[33]}});
    result = result | (input_34 & {2{sel[34]}});
    result = result | (input_35 & {2{sel[35]}});
    result = result | (input_36 & {2{sel[36]}});
    result = result | (input_37 & {2{sel[37]}});
    result = result | (input_38 & {2{sel[38]}});
    result = result | (input_39 & {2{sel[39]}});
    result = result | (input_40 & {2{sel[40]}});
    result = result | (input_41 & {2{sel[41]}});
    result = result | (input_42 & {2{sel[42]}});
    result = result | (input_43 & {2{sel[43]}});
    result = result | (input_44 & {2{sel[44]}});
    result = result | (input_45 & {2{sel[45]}});
    result = result | (input_46 & {2{sel[46]}});
    result = result | (input_47 & {2{sel[47]}});
    result = result | (input_48 & {2{sel[48]}});
    result = result | (input_49 & {2{sel[49]}});
    result = result | (input_50 & {2{sel[50]}});
    MUX1HOT_v_2_51_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_32_2;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [31:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    MUX1HOT_v_4_32_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_34_2;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [33:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    MUX1HOT_v_4_34_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_35_2;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [34:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    MUX1HOT_v_4_35_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_49_2;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [48:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    MUX1HOT_v_4_49_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_51_2;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [50:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    MUX1HOT_v_4_51_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_65_2;
    input [4:0] input_64;
    input [4:0] input_63;
    input [4:0] input_62;
    input [4:0] input_61;
    input [4:0] input_60;
    input [4:0] input_59;
    input [4:0] input_58;
    input [4:0] input_57;
    input [4:0] input_56;
    input [4:0] input_55;
    input [4:0] input_54;
    input [4:0] input_53;
    input [4:0] input_52;
    input [4:0] input_51;
    input [4:0] input_50;
    input [4:0] input_49;
    input [4:0] input_48;
    input [4:0] input_47;
    input [4:0] input_46;
    input [4:0] input_45;
    input [4:0] input_44;
    input [4:0] input_43;
    input [4:0] input_42;
    input [4:0] input_41;
    input [4:0] input_40;
    input [4:0] input_39;
    input [4:0] input_38;
    input [4:0] input_37;
    input [4:0] input_36;
    input [4:0] input_35;
    input [4:0] input_34;
    input [4:0] input_33;
    input [4:0] input_32;
    input [4:0] input_31;
    input [4:0] input_30;
    input [4:0] input_29;
    input [4:0] input_28;
    input [4:0] input_27;
    input [4:0] input_26;
    input [4:0] input_25;
    input [4:0] input_24;
    input [4:0] input_23;
    input [4:0] input_22;
    input [4:0] input_21;
    input [4:0] input_20;
    input [4:0] input_19;
    input [4:0] input_18;
    input [4:0] input_17;
    input [4:0] input_16;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [64:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    result = result | (input_13 & {5{sel[13]}});
    result = result | (input_14 & {5{sel[14]}});
    result = result | (input_15 & {5{sel[15]}});
    result = result | (input_16 & {5{sel[16]}});
    result = result | (input_17 & {5{sel[17]}});
    result = result | (input_18 & {5{sel[18]}});
    result = result | (input_19 & {5{sel[19]}});
    result = result | (input_20 & {5{sel[20]}});
    result = result | (input_21 & {5{sel[21]}});
    result = result | (input_22 & {5{sel[22]}});
    result = result | (input_23 & {5{sel[23]}});
    result = result | (input_24 & {5{sel[24]}});
    result = result | (input_25 & {5{sel[25]}});
    result = result | (input_26 & {5{sel[26]}});
    result = result | (input_27 & {5{sel[27]}});
    result = result | (input_28 & {5{sel[28]}});
    result = result | (input_29 & {5{sel[29]}});
    result = result | (input_30 & {5{sel[30]}});
    result = result | (input_31 & {5{sel[31]}});
    result = result | (input_32 & {5{sel[32]}});
    result = result | (input_33 & {5{sel[33]}});
    result = result | (input_34 & {5{sel[34]}});
    result = result | (input_35 & {5{sel[35]}});
    result = result | (input_36 & {5{sel[36]}});
    result = result | (input_37 & {5{sel[37]}});
    result = result | (input_38 & {5{sel[38]}});
    result = result | (input_39 & {5{sel[39]}});
    result = result | (input_40 & {5{sel[40]}});
    result = result | (input_41 & {5{sel[41]}});
    result = result | (input_42 & {5{sel[42]}});
    result = result | (input_43 & {5{sel[43]}});
    result = result | (input_44 & {5{sel[44]}});
    result = result | (input_45 & {5{sel[45]}});
    result = result | (input_46 & {5{sel[46]}});
    result = result | (input_47 & {5{sel[47]}});
    result = result | (input_48 & {5{sel[48]}});
    result = result | (input_49 & {5{sel[49]}});
    result = result | (input_50 & {5{sel[50]}});
    result = result | (input_51 & {5{sel[51]}});
    result = result | (input_52 & {5{sel[52]}});
    result = result | (input_53 & {5{sel[53]}});
    result = result | (input_54 & {5{sel[54]}});
    result = result | (input_55 & {5{sel[55]}});
    result = result | (input_56 & {5{sel[56]}});
    result = result | (input_57 & {5{sel[57]}});
    result = result | (input_58 & {5{sel[58]}});
    result = result | (input_59 & {5{sel[59]}});
    result = result | (input_60 & {5{sel[60]}});
    result = result | (input_61 & {5{sel[61]}});
    result = result | (input_62 & {5{sel[62]}});
    result = result | (input_63 & {5{sel[63]}});
    result = result | (input_64 & {5{sel[64]}});
    MUX1HOT_v_5_65_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_5_2;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [4:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    MUX1HOT_v_7_5_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [4:0] signext_5_4;
    input [3:0] vector;
  begin
    signext_5_4= {{1{vector[3]}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_4;
    input [3:0] vector;
  begin
    signext_7_4= {{3{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [7:0] conv_s2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_4_7 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_7 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_m_rsc_dat, input_m_triosy_lz, input_e_rsc_dat, input_e_triosy_lz,
      taps_m_rsc_dat, taps_m_triosy_lz, taps_e_rsc_dat, taps_e_triosy_lz, return_m_rsc_dat,
      return_m_triosy_lz, return_e_rsc_dat, return_e_triosy_lz
);
  input clk;
  input rst;
  input [10:0] input_m_rsc_dat;
  output input_m_triosy_lz;
  input [4:0] input_e_rsc_dat;
  output input_e_triosy_lz;
  input [351:0] taps_m_rsc_dat;
  output taps_m_triosy_lz;
  input [159:0] taps_e_rsc_dat;
  output taps_e_triosy_lz;
  output [10:0] return_m_rsc_dat;
  output return_m_triosy_lz;
  output [4:0] return_e_rsc_dat;
  output return_e_triosy_lz;


  // Interconnect Declarations
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;


  // Interconnect Declarations for Component Instantiations 
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_1 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_2 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_3 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_4 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_5 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_6 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_7 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_8 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_9 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_10 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_11 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_12 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_13 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_14 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_15 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_16 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_17 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_18 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_19 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_20 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_21 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_22 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_23 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_24 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_25 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_26 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_27 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_28 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_29 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_30 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_31 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn)
    );
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .input_m_rsc_dat(input_m_rsc_dat),
      .input_m_triosy_lz(input_m_triosy_lz),
      .input_e_rsc_dat(input_e_rsc_dat),
      .input_e_triosy_lz(input_e_triosy_lz),
      .taps_m_rsc_dat(taps_m_rsc_dat),
      .taps_m_triosy_lz(taps_m_triosy_lz),
      .taps_e_rsc_dat(taps_e_rsc_dat),
      .taps_e_triosy_lz(taps_e_triosy_lz),
      .return_m_rsc_dat(return_m_rsc_dat),
      .return_m_triosy_lz(return_m_triosy_lz),
      .return_e_rsc_dat(return_e_rsc_dat),
      .return_e_triosy_lz(return_e_triosy_lz),
      .MAC_1_leading_sign_18_1_1_0_cmp_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn)
    );
endmodule



