
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v5.v 
module mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/leading_sign_13_1_1_0_fbd6b6484e0226fdfa7c7e6838ce99f45fe9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:36 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_13_1_1_0
// ------------------------------------------------------------------


module leading_sign_13_1_1_0 (
  mantissa, all_same, rtn
);
  input [12:0] mantissa;
  output all_same;
  output [3:0] rtn;


  // Interconnect Declarations
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire [11:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0;
  wire c_h_1_2;
  wire c_h_1_4;

  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0 = (mantissa[11:0])
      ^ (signext_12_1(~ (mantissa[12])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[9:8]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11:10]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7:6]==2'b11);
  assign c_h_1_2 = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[5:4]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3:2]==2'b11);
  assign c_h_1_4 = c_h_1_2 & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[1:0]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1 &
      c_h_1_4;
  assign all_same = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      = (c_h_1_2 & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3))
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl = ~(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      | (~ c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl = ~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[10:9]!=2'b10))
      & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[6:5]!=2'b10))))
      & c_h_1_2)) & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[2:1]!=2'b10))))
      & c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl
      = ~(MUX_v_2_2_2(({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl}), 2'b11,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4));
  assign rtn = {c_h_1_4 , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl};

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [11:0] signext_12_1;
    input  vector;
  begin
    signext_12_1= {{11{vector}}, vector};
  end
  endfunction

endmodule




//------> ../td_ccore_solutions/leading_sign_18_1_1_0_7b2153b3b691fe1ab68d43c72c494a7b6845_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:37 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_18_1_1_0
// ------------------------------------------------------------------


module leading_sign_18_1_1_0 (
  mantissa, all_same, rtn
);
  input [17:0] mantissa;
  output all_same;
  output [4:0] rtn;


  // Interconnect Declarations
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1;
  wire [16:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_7;

  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0
      = (mantissa[16:0]) ^ (signext_17_1(~ (mantissa[17])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[14:13]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16:15]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12:11]==2'b11);
  assign c_h_1_2 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[10:9]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[6:5]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8:7]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4:3]==2'b11);
  assign c_h_1_5 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[2:1]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[0])
      & c_h_1_7;
  assign all_same = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      = c_h_1_6 & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3))
      & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl
      = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[15:14]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[11:10]!=2'b10))))
      & c_h_1_2)) & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[7:6]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[3:2]!=2'b10))))
      & c_h_1_5)))) & c_h_1_6)) & (~ c_h_1_7)) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign rtn = {c_h_1_7 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl};

  function automatic [16:0] signext_17_1;
    input  vector;
  begin
    signext_17_1= {{16{vector}}, vector};
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Wed Apr 23 23:11:12 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [6:0] fsm_output;
  reg [6:0] fsm_output;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 7'd0,
    main_C_1 = 7'd1,
    main_C_2 = 7'd2,
    main_C_3 = 7'd3,
    main_C_4 = 7'd4,
    main_C_5 = 7'd5,
    main_C_6 = 7'd6,
    main_C_7 = 7'd7,
    main_C_8 = 7'd8,
    main_C_9 = 7'd9,
    main_C_10 = 7'd10,
    main_C_11 = 7'd11,
    main_C_12 = 7'd12,
    main_C_13 = 7'd13,
    main_C_14 = 7'd14,
    main_C_15 = 7'd15,
    main_C_16 = 7'd16,
    main_C_17 = 7'd17,
    main_C_18 = 7'd18,
    main_C_19 = 7'd19,
    main_C_20 = 7'd20,
    main_C_21 = 7'd21,
    main_C_22 = 7'd22,
    main_C_23 = 7'd23,
    main_C_24 = 7'd24,
    main_C_25 = 7'd25,
    main_C_26 = 7'd26,
    main_C_27 = 7'd27,
    main_C_28 = 7'd28,
    main_C_29 = 7'd29,
    main_C_30 = 7'd30,
    main_C_31 = 7'd31,
    main_C_32 = 7'd32,
    main_C_33 = 7'd33,
    main_C_34 = 7'd34,
    main_C_35 = 7'd35,
    main_C_36 = 7'd36,
    main_C_37 = 7'd37,
    main_C_38 = 7'd38,
    main_C_39 = 7'd39,
    main_C_40 = 7'd40,
    main_C_41 = 7'd41,
    main_C_42 = 7'd42,
    main_C_43 = 7'd43,
    main_C_44 = 7'd44,
    main_C_45 = 7'd45,
    main_C_46 = 7'd46,
    main_C_47 = 7'd47,
    main_C_48 = 7'd48,
    main_C_49 = 7'd49,
    main_C_50 = 7'd50,
    main_C_51 = 7'd51,
    main_C_52 = 7'd52,
    main_C_53 = 7'd53,
    main_C_54 = 7'd54,
    main_C_55 = 7'd55,
    main_C_56 = 7'd56,
    main_C_57 = 7'd57,
    main_C_58 = 7'd58,
    main_C_59 = 7'd59,
    main_C_60 = 7'd60,
    main_C_61 = 7'd61,
    main_C_62 = 7'd62,
    main_C_63 = 7'd63,
    main_C_64 = 7'd64,
    main_C_65 = 7'd65,
    main_C_66 = 7'd66,
    main_C_67 = 7'd67,
    main_C_68 = 7'd68,
    main_C_69 = 7'd69,
    main_C_70 = 7'd70;

  reg [6:0] state_var;
  reg [6:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 7'b0000001;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 7'b0000010;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 7'b0000011;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 7'b0000100;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 7'b0000101;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 7'b0000110;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 7'b0000111;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 7'b0001000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 7'b0001001;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 7'b0001010;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 7'b0001011;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 7'b0001100;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 7'b0001101;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 7'b0001110;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 7'b0001111;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 7'b0010000;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 7'b0010001;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 7'b0010010;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 7'b0010011;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 7'b0010100;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 7'b0010101;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 7'b0010110;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 7'b0010111;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 7'b0011000;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 7'b0011001;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 7'b0011010;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 7'b0011011;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 7'b0011100;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 7'b0011101;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 7'b0011110;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 7'b0011111;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 7'b0100000;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 7'b0100001;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 7'b0100010;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 7'b0100011;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 7'b0100100;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 7'b0100101;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 7'b0100110;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 7'b0100111;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 7'b0101000;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 7'b0101001;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 7'b0101010;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 7'b0101011;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 7'b0101100;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 7'b0101101;
        state_var_NS = main_C_46;
      end
      main_C_46 : begin
        fsm_output = 7'b0101110;
        state_var_NS = main_C_47;
      end
      main_C_47 : begin
        fsm_output = 7'b0101111;
        state_var_NS = main_C_48;
      end
      main_C_48 : begin
        fsm_output = 7'b0110000;
        state_var_NS = main_C_49;
      end
      main_C_49 : begin
        fsm_output = 7'b0110001;
        state_var_NS = main_C_50;
      end
      main_C_50 : begin
        fsm_output = 7'b0110010;
        state_var_NS = main_C_51;
      end
      main_C_51 : begin
        fsm_output = 7'b0110011;
        state_var_NS = main_C_52;
      end
      main_C_52 : begin
        fsm_output = 7'b0110100;
        state_var_NS = main_C_53;
      end
      main_C_53 : begin
        fsm_output = 7'b0110101;
        state_var_NS = main_C_54;
      end
      main_C_54 : begin
        fsm_output = 7'b0110110;
        state_var_NS = main_C_55;
      end
      main_C_55 : begin
        fsm_output = 7'b0110111;
        state_var_NS = main_C_56;
      end
      main_C_56 : begin
        fsm_output = 7'b0111000;
        state_var_NS = main_C_57;
      end
      main_C_57 : begin
        fsm_output = 7'b0111001;
        state_var_NS = main_C_58;
      end
      main_C_58 : begin
        fsm_output = 7'b0111010;
        state_var_NS = main_C_59;
      end
      main_C_59 : begin
        fsm_output = 7'b0111011;
        state_var_NS = main_C_60;
      end
      main_C_60 : begin
        fsm_output = 7'b0111100;
        state_var_NS = main_C_61;
      end
      main_C_61 : begin
        fsm_output = 7'b0111101;
        state_var_NS = main_C_62;
      end
      main_C_62 : begin
        fsm_output = 7'b0111110;
        state_var_NS = main_C_63;
      end
      main_C_63 : begin
        fsm_output = 7'b0111111;
        state_var_NS = main_C_64;
      end
      main_C_64 : begin
        fsm_output = 7'b1000000;
        state_var_NS = main_C_65;
      end
      main_C_65 : begin
        fsm_output = 7'b1000001;
        state_var_NS = main_C_66;
      end
      main_C_66 : begin
        fsm_output = 7'b1000010;
        state_var_NS = main_C_67;
      end
      main_C_67 : begin
        fsm_output = 7'b1000011;
        state_var_NS = main_C_68;
      end
      main_C_68 : begin
        fsm_output = 7'b1000100;
        state_var_NS = main_C_69;
      end
      main_C_69 : begin
        fsm_output = 7'b1000101;
        state_var_NS = main_C_70;
      end
      main_C_70 : begin
        fsm_output = 7'b1000110;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 7'b0000000;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core_wait_dp
// ------------------------------------------------------------------


module fir_core_wait_dp (
  clk, rst, MAC_1_leading_sign_18_1_1_0_cmp_all_same, MAC_1_leading_sign_18_1_1_0_cmp_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same, MAC_1_leading_sign_18_1_1_0_cmp_32_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same, MAC_1_leading_sign_18_1_1_0_cmp_33_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same, MAC_1_leading_sign_18_1_1_0_cmp_34_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same, MAC_1_leading_sign_18_1_1_0_cmp_35_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same, MAC_1_leading_sign_18_1_1_0_cmp_36_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same, MAC_1_leading_sign_18_1_1_0_cmp_37_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same, MAC_1_leading_sign_18_1_1_0_cmp_38_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same, MAC_1_leading_sign_18_1_1_0_cmp_39_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same, MAC_1_leading_sign_18_1_1_0_cmp_40_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same, MAC_1_leading_sign_18_1_1_0_cmp_41_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same, MAC_1_leading_sign_18_1_1_0_cmp_42_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same, MAC_1_leading_sign_18_1_1_0_cmp_43_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same, MAC_1_leading_sign_18_1_1_0_cmp_44_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same, MAC_1_leading_sign_18_1_1_0_cmp_45_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same, MAC_1_leading_sign_18_1_1_0_cmp_46_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same, MAC_1_leading_sign_18_1_1_0_cmp_47_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same, MAC_1_leading_sign_18_1_1_0_cmp_48_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same, MAC_1_leading_sign_18_1_1_0_cmp_49_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same, MAC_1_leading_sign_18_1_1_0_cmp_50_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same, MAC_1_leading_sign_18_1_1_0_cmp_51_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same, MAC_1_leading_sign_18_1_1_0_cmp_52_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same, MAC_1_leading_sign_18_1_1_0_cmp_53_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same, MAC_1_leading_sign_18_1_1_0_cmp_54_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same, MAC_1_leading_sign_18_1_1_0_cmp_55_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same, MAC_1_leading_sign_18_1_1_0_cmp_56_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same, MAC_1_leading_sign_18_1_1_0_cmp_57_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same, MAC_1_leading_sign_18_1_1_0_cmp_58_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same, MAC_1_leading_sign_18_1_1_0_cmp_59_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same, MAC_1_leading_sign_18_1_1_0_cmp_60_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same, MAC_1_leading_sign_18_1_1_0_cmp_61_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same, MAC_1_leading_sign_18_1_1_0_cmp_62_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same, MAC_1_leading_sign_18_1_1_0_cmp_63_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg
);
  input clk;
  input rst;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;
  output MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;


  // Interconnect Declarations
  reg MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg;


  // Interconnect Declarations for Component Instantiations 
  assign MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg;
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg <= 5'b00000;
    end
    else begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, input_real_m_rsc_dat, input_real_m_triosy_lz, input_real_e_rsc_dat, input_real_e_triosy_lz,
      input_imag_m_rsc_dat, input_imag_m_triosy_lz, input_imag_e_rsc_dat, input_imag_e_triosy_lz,
      taps_real_m_rsc_dat, taps_real_m_triosy_lz, taps_real_e_rsc_dat, taps_real_e_triosy_lz,
      taps_imag_m_rsc_dat, taps_imag_m_triosy_lz, taps_imag_e_rsc_dat, taps_imag_e_triosy_lz,
      return_real_m_rsc_dat, return_real_m_triosy_lz, return_real_e_rsc_dat, return_real_e_triosy_lz,
      return_imag_m_rsc_dat, return_imag_m_triosy_lz, return_imag_e_rsc_dat, return_imag_e_triosy_lz,
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_rtn, MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_2_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn, MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_4_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn, MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_6_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn, MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_8_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn, MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_10_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn, MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_12_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn, MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_14_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn, MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_16_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn, MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_18_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn, MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_20_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn, MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_22_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn, MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_24_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn, MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_26_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn, MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_28_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn, MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_30_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn, MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_32_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_32_rtn, MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same, MAC_1_leading_sign_18_1_1_0_cmp_33_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_34_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_34_rtn, MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same, MAC_1_leading_sign_18_1_1_0_cmp_35_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_36_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_36_rtn, MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same, MAC_1_leading_sign_18_1_1_0_cmp_37_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_38_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_38_rtn, MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same, MAC_1_leading_sign_18_1_1_0_cmp_39_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_40_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_40_rtn, MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same, MAC_1_leading_sign_18_1_1_0_cmp_41_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_42_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_42_rtn, MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same, MAC_1_leading_sign_18_1_1_0_cmp_43_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_44_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_44_rtn, MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same, MAC_1_leading_sign_18_1_1_0_cmp_45_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_46_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_46_rtn, MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same, MAC_1_leading_sign_18_1_1_0_cmp_47_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_48_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_48_rtn, MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same, MAC_1_leading_sign_18_1_1_0_cmp_49_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_50_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_50_rtn, MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same, MAC_1_leading_sign_18_1_1_0_cmp_51_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_52_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_52_rtn, MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same, MAC_1_leading_sign_18_1_1_0_cmp_53_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_54_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_54_rtn, MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same, MAC_1_leading_sign_18_1_1_0_cmp_55_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_56_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_56_rtn, MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same, MAC_1_leading_sign_18_1_1_0_cmp_57_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_58_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_58_rtn, MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same, MAC_1_leading_sign_18_1_1_0_cmp_59_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_60_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_60_rtn, MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same, MAC_1_leading_sign_18_1_1_0_cmp_61_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_62_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_62_rtn, MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same, MAC_1_leading_sign_18_1_1_0_cmp_63_rtn
);
  input clk;
  input rst;
  input [10:0] input_real_m_rsc_dat;
  output input_real_m_triosy_lz;
  input [4:0] input_real_e_rsc_dat;
  output input_real_e_triosy_lz;
  input [10:0] input_imag_m_rsc_dat;
  output input_imag_m_triosy_lz;
  input [4:0] input_imag_e_rsc_dat;
  output input_imag_e_triosy_lz;
  input [175:0] taps_real_m_rsc_dat;
  output taps_real_m_triosy_lz;
  input [79:0] taps_real_e_rsc_dat;
  output taps_real_e_triosy_lz;
  input [175:0] taps_imag_m_rsc_dat;
  output taps_imag_m_triosy_lz;
  input [79:0] taps_imag_e_rsc_dat;
  output taps_imag_e_triosy_lz;
  output [10:0] return_real_m_rsc_dat;
  output return_real_m_triosy_lz;
  output [4:0] return_real_e_rsc_dat;
  output return_real_e_triosy_lz;
  output [10:0] return_imag_m_rsc_dat;
  output return_imag_m_triosy_lz;
  output [4:0] return_imag_e_rsc_dat;
  output return_imag_e_triosy_lz;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;


  // Interconnect Declarations
  wire [10:0] input_real_m_rsci_idat;
  wire [4:0] input_real_e_rsci_idat;
  wire [10:0] input_imag_m_rsci_idat;
  wire [4:0] input_imag_e_rsci_idat;
  wire [175:0] taps_real_m_rsci_idat;
  wire [79:0] taps_real_e_rsci_idat;
  wire [175:0] taps_imag_m_rsci_idat;
  wire [79:0] taps_imag_e_rsci_idat;
  reg [10:0] return_real_m_rsci_idat;
  reg [4:0] return_real_e_rsci_idat;
  reg [10:0] return_imag_m_rsci_idat;
  reg [4:0] return_imag_e_rsci_idat;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;
  wire [6:0] fsm_output;
  wire [5:0] MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp;
  wire [5:0] MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp;
  wire [5:0] MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp;
  wire MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp;
  wire [5:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [5:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [5:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [5:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [5:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_12_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_11_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_10_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_10_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_10_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_10_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [5:0] MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp;
  wire [5:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_16_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp;
  wire [5:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_15_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_16_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp;
  wire [5:0] MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_8_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_8_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_8_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_7_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_7_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_7_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_6_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_6_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_6_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_5_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_5_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_5_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_4_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_4_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_4_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_3_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_3_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_3_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_2_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_2_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_2_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [5:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire [6:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp;
  wire MAC_1_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  wire MAC_1_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  wire [5:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_1_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  wire MAC_1_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  wire [2:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire and_dcpl_2;
  wire or_tmp_20;
  wire mux_tmp_31;
  wire mux_tmp_56;
  wire nor_tmp_6;
  wire not_tmp_212;
  wire mux_tmp_65;
  wire or_dcpl_193;
  wire or_dcpl_194;
  wire or_dcpl_195;
  wire or_dcpl_196;
  wire or_dcpl_197;
  wire and_dcpl_164;
  wire and_dcpl_166;
  wire and_dcpl_167;
  wire and_dcpl_169;
  wire or_dcpl_200;
  wire or_dcpl_201;
  wire or_dcpl_204;
  wire and_dcpl_182;
  wire and_dcpl_183;
  wire and_dcpl_184;
  wire and_dcpl_185;
  wire and_dcpl_186;
  wire and_dcpl_187;
  wire and_dcpl_188;
  wire and_dcpl_189;
  wire or_dcpl_207;
  wire and_dcpl_190;
  wire and_dcpl_191;
  wire and_dcpl_192;
  wire and_dcpl_193;
  wire and_dcpl_194;
  wire and_dcpl_195;
  wire and_dcpl_196;
  wire and_dcpl_197;
  wire and_dcpl_198;
  wire and_dcpl_199;
  wire and_dcpl_200;
  wire xor_dcpl;
  wire and_dcpl_202;
  wire and_dcpl_203;
  wire and_dcpl_206;
  wire and_dcpl_208;
  wire and_dcpl_209;
  wire and_dcpl_210;
  wire and_dcpl_211;
  wire and_dcpl_212;
  wire or_tmp_98;
  wire or_tmp_100;
  wire mux_tmp_98;
  wire mux_tmp_99;
  wire and_dcpl_213;
  wire or_tmp_102;
  wire mux_tmp_101;
  wire or_tmp_104;
  wire and_dcpl_215;
  wire and_dcpl_218;
  wire or_tmp_107;
  wire and_dcpl_220;
  wire and_dcpl_222;
  wire and_dcpl_223;
  wire or_tmp_111;
  wire mux_tmp_121;
  wire and_dcpl_227;
  wire and_dcpl_231;
  wire and_dcpl_232;
  wire mux_tmp_143;
  wire and_dcpl_243;
  wire mux_tmp_146;
  wire mux_tmp_147;
  wire mux_tmp_149;
  wire mux_tmp_150;
  wire not_tmp_284;
  wire and_dcpl_245;
  wire and_dcpl_248;
  wire and_dcpl_251;
  wire and_dcpl_254;
  wire and_dcpl_257;
  wire or_tmp_131;
  wire and_dcpl_260;
  wire and_dcpl_277;
  wire and_dcpl_280;
  wire and_dcpl_281;
  wire and_dcpl_282;
  wire and_dcpl_283;
  wire and_dcpl_284;
  wire and_dcpl_285;
  wire and_dcpl_286;
  wire and_dcpl_287;
  wire and_dcpl_288;
  wire and_dcpl_289;
  wire and_dcpl_290;
  wire and_dcpl_291;
  wire and_dcpl_292;
  wire and_dcpl_293;
  wire and_dcpl_294;
  wire and_dcpl_295;
  wire and_dcpl_296;
  wire and_dcpl_297;
  wire and_dcpl_298;
  wire and_dcpl_299;
  wire and_dcpl_300;
  wire and_dcpl_327;
  wire and_dcpl_345;
  wire mux_tmp_188;
  wire not_tmp_307;
  wire mux_tmp_223;
  wire or_dcpl_229;
  wire and_dcpl_361;
  wire and_dcpl_364;
  wire and_dcpl_367;
  wire and_dcpl_370;
  wire and_dcpl_373;
  wire and_dcpl_376;
  wire and_dcpl_379;
  wire and_dcpl_382;
  wire and_dcpl_385;
  wire and_dcpl_388;
  wire and_dcpl_392;
  wire and_dcpl_395;
  wire and_dcpl_399;
  wire and_dcpl_402;
  wire and_dcpl_405;
  wire and_dcpl_408;
  wire and_dcpl_409;
  wire mux_tmp_236;
  wire and_dcpl_420;
  wire and_dcpl_423;
  wire and_dcpl_426;
  wire and_dcpl_429;
  wire and_dcpl_432;
  wire and_dcpl_435;
  wire and_dcpl_452;
  wire and_dcpl_455;
  wire or_tmp_153;
  wire or_tmp_154;
  wire and_dcpl_478;
  wire and_dcpl_481;
  wire and_dcpl_482;
  wire and_dcpl_484;
  wire and_dcpl_485;
  wire and_dcpl_487;
  wire and_dcpl_496;
  wire and_dcpl_499;
  wire and_dcpl_521;
  wire and_dcpl_524;
  wire nor_tmp_26;
  wire mux_tmp_247;
  wire and_dcpl_552;
  wire and_dcpl_555;
  wire and_dcpl_574;
  wire mux_tmp_257;
  wire and_dcpl_596;
  wire and_dcpl_599;
  wire mux_tmp_261;
  wire and_dcpl_624;
  wire and_dcpl_633;
  wire nor_tmp_29;
  wire and_dcpl_637;
  wire and_dcpl_640;
  wire and_dcpl_647;
  wire and_dcpl_654;
  wire and_dcpl_655;
  wire and_dcpl_663;
  wire and_dcpl_669;
  wire and_dcpl_679;
  wire and_dcpl_689;
  wire and_dcpl_692;
  wire and_dcpl_720;
  wire and_dcpl_723;
  wire and_dcpl_799;
  wire and_dcpl_802;
  wire and_dcpl_854;
  wire and_dcpl_857;
  wire and_dcpl_937;
  wire and_dcpl_963;
  wire and_dcpl_964;
  wire and_dcpl_976;
  wire and_dcpl_981;
  wire and_dcpl_985;
  wire and_dcpl_990;
  wire or_dcpl_257;
  wire or_tmp_238;
  wire and_dcpl_1012;
  wire or_dcpl_262;
  wire and_dcpl_1017;
  wire and_dcpl_1036;
  wire and_dcpl_1054;
  wire and_dcpl_1070;
  wire and_dcpl_1077;
  wire and_dcpl_1078;
  wire and_dcpl_1082;
  wire and_dcpl_1090;
  wire and_dcpl_1097;
  wire and_dcpl_1098;
  wire and_dcpl_1102;
  wire and_dcpl_1106;
  wire and_dcpl_1110;
  wire and_dcpl_1138;
  wire and_dcpl_1142;
  wire and_dcpl_1173;
  wire and_dcpl_1187;
  wire and_dcpl_1218;
  wire mux_tmp_380;
  wire and_dcpl_1267;
  wire mux_tmp_384;
  wire mux_tmp_393;
  wire or_tmp_275;
  wire mux_tmp_402;
  wire and_dcpl_1355;
  wire or_tmp_291;
  wire and_dcpl_1363;
  wire and_dcpl_1366;
  wire and_dcpl_1369;
  wire and_dcpl_1374;
  wire or_tmp_300;
  wire or_tmp_303;
  wire and_dcpl_1383;
  wire and_dcpl_1389;
  wire and_dcpl_1395;
  wire and_dcpl_1398;
  wire or_tmp_319;
  wire not_tmp_606;
  wire and_dcpl_1413;
  wire and_dcpl_1425;
  wire and_dcpl_1426;
  wire and_dcpl_1427;
  wire and_dcpl_1428;
  wire and_dcpl_1429;
  wire and_dcpl_1430;
  wire and_dcpl_1431;
  wire and_dcpl_1432;
  wire and_dcpl_1433;
  wire and_dcpl_1434;
  wire and_dcpl_1435;
  wire and_dcpl_1436;
  wire and_dcpl_1437;
  wire and_dcpl_1438;
  wire and_dcpl_1439;
  wire and_dcpl_1440;
  wire and_dcpl_1450;
  wire and_dcpl_1463;
  wire mux_tmp_477;
  wire mux_tmp_481;
  wire mux_tmp_483;
  wire and_dcpl_1547;
  wire and_dcpl_1550;
  wire and_dcpl_1551;
  wire and_dcpl_1554;
  wire and_dcpl_1557;
  wire and_dcpl_1562;
  wire and_dcpl_1565;
  wire and_dcpl_1568;
  wire and_dcpl_1575;
  wire and_dcpl_1578;
  wire or_dcpl_485;
  wire or_dcpl_486;
  wire or_dcpl_507;
  wire or_dcpl_509;
  wire and_dcpl_1579;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6;
  reg MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm;
  reg ac_float_cctor_operator_return_59_sva;
  reg MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_32_sva;
  reg MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_operator_return_31_sva;
  reg MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_30_sva;
  reg MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_operator_return_3_sva;
  reg MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_48_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm;
  reg ac_float_cctor_operator_return_42_sva;
  reg MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_operator_return_17_sva;
  reg MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_12_sva;
  reg MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_operator_return_63_sva;
  reg MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_62_sva;
  reg MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_61_sva;
  reg MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_operator_return_60_sva;
  reg MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_operator_return_29_sva;
  reg MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm;
  wire [10:0] operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_15_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_14_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva;
  wire [10:0] operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_14_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  wire [10:0] operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_13_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva;
  wire [10:0] operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_13_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  wire [10:0] operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_12_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva;
  wire [10:0] operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_12_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  wire [10:0] operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_11_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva;
  wire [10:0] operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_11_lpi_1_dfm_1;
  reg MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva;
  reg MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  wire [10:0] operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1;
  wire [10:0] operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_9_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_8_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_9_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm;
  wire [10:0] operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2;
  wire [10:0] operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_9_lpi_1_dfm_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva;
  reg MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva;
  reg MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva;
  reg MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva;
  reg MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  reg [10:0] delay_lane_imag_m_14_sva;
  reg [10:0] delay_lane_real_m_14_sva;
  reg [10:0] delay_lane_imag_m_13_sva;
  reg [10:0] delay_lane_real_m_13_sva;
  reg [10:0] delay_lane_imag_m_12_sva;
  reg [10:0] delay_lane_real_m_12_sva;
  reg [10:0] delay_lane_imag_m_11_sva;
  reg [10:0] delay_lane_real_m_11_sva;
  reg [10:0] delay_lane_imag_m_10_sva;
  reg [10:0] delay_lane_real_m_10_sva;
  reg [10:0] delay_lane_imag_m_9_sva;
  reg [10:0] delay_lane_real_m_9_sva;
  reg [10:0] delay_lane_imag_m_8_sva;
  reg [10:0] delay_lane_real_m_8_sva;
  reg [10:0] delay_lane_imag_m_7_sva;
  reg [10:0] delay_lane_real_m_7_sva;
  reg [10:0] delay_lane_imag_m_6_sva;
  reg [10:0] delay_lane_real_m_6_sva;
  reg [10:0] delay_lane_imag_m_5_sva;
  reg [10:0] delay_lane_real_m_5_sva;
  reg [10:0] delay_lane_imag_m_4_sva;
  reg [10:0] delay_lane_real_m_4_sva;
  reg [10:0] delay_lane_imag_m_3_sva;
  reg [10:0] delay_lane_real_m_3_sva;
  reg [10:0] delay_lane_imag_m_2_sva;
  reg [10:0] delay_lane_real_m_2_sva;
  reg [10:0] delay_lane_imag_m_1_sva;
  reg [10:0] delay_lane_real_m_1_sva;
  reg [10:0] delay_lane_imag_m_0_sva;
  reg [10:0] delay_lane_real_m_0_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1;
  wire [4:0] operator_i_e_1_lpi_1_dfm_mx0;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_22;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_26;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_38;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_40;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_42;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_19;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_28;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_32;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_16;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_36;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_17;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_18;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva;
  reg [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva;
  wire ac_float_cctor_operator_return_2_sva_mx0w2;
  wire ac_float_cctor_operator_return_48_sva_mx0w2;
  wire ac_float_cctor_operator_return_47_sva_mx0w2;
  wire ac_float_cctor_operator_return_17_sva_mx0w2;
  wire ac_float_cctor_operator_return_46_sva_mx0w2;
  wire ac_float_cctor_operator_return_16_sva_mx0w2;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_15_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_14_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_14_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_13_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_13_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_12_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_12_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_11_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_11_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1;
  wire ac_float_cctor_operator_return_42_sva_mx0w1;
  wire ac_float_cctor_operator_return_57_sva_mx0w1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_9_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_9_lpi_1_dfm_mx0;
  wire ac_float_cctor_operator_return_12_sva_mx0w1;
  wire ac_float_cctor_operator_return_27_sva_mx0w1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_9_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
  reg [4:0] operator_ac_float_cctor_e_29_lpi_1_dfm;
  reg [4:0] operator_ac_float_cctor_e_19_lpi_1_dfm;
  reg [4:0] operator_ac_float_cctor_e_14_lpi_1_dfm;
  reg [4:0] operator_ac_float_cctor_e_65_lpi_1_dfm;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva;
  reg [4:0] operator_ac_float_cctor_e_64_lpi_1_dfm;
  reg [4:0] operator_ac_float_cctor_e_3_lpi_1_dfm;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva;
  wire [6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_seb;
  wire and_362_ssc;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1;
  wire [11:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt;
  wire [12:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7;
  wire [11:0] MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt;
  wire [12:0] nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_1_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_11_7;
  wire [11:0] MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_1_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_11_7;
  wire [11:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_8_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7;
  wire and_1501_m1c;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0;
  wire [11:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_4_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_11;
  wire [11:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_3_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_11;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_2_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_11;
  wire [11:0] MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_5_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_11;
  wire [11:0] MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_7_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_11;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_6_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_11;
  reg [3:0] MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0;
  reg [3:0] MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_or_cse;
  reg reg_return_imag_e_triosy_obj_ld_cse;
  reg reg_taps_imag_e_triosy_obj_ld_cse;
  wire or_6_cse;
  wire nor_478_cse;
  wire nor_81_cse;
  wire or_972_cse;
  wire or_467_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_2_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_1_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_3_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_1_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_4_cse;
  wire and_1628_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_8_cse;
  wire nor_522_cse;
  wire nor_521_cse;
  wire nor_524_cse;
  wire nor_523_cse;
  wire nor_540_cse;
  wire nor_539_cse;
  wire nor_542_cse;
  wire nor_541_cse;
  wire [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse;
  wire nor_137_cse;
  wire or_361_cse;
  wire nor_469_cse;
  wire nor_98_cse;
  wire and_1593_cse;
  wire or_966_cse;
  wire or_730_cse;
  wire or_967_cse;
  wire or_968_cse;
  wire nor_195_cse;
  wire nor_199_cse;
  wire or_900_cse;
  wire nor_479_cse;
  wire nor_75_cse;
  wire nor_429_cse;
  wire nor_200_cse;
  wire nor_442_cse;
  wire nor_450_cse;
  wire nor_56_cse;
  wire nor_203_cse;
  wire nor_456_cse;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_ssc;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_11_7;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_5_ssc;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_11_7;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_11_7;
  wire [4:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  wire [4:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [4:0] MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  wire [4:0] MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  wire [4:0] MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  wire [4:0] MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb;
  wire [4:0] MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb;
  wire [4:0] MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb;
  wire [4:0] MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb;
  wire [4:0] MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb;
  wire [4:0] MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb;
  wire [4:0] MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb;
  wire [4:0] MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb;
  wire [4:0] MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb;
  wire [4:0] MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb;
  wire [4:0] MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb;
  wire [4:0] MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb;
  reg MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4;
  reg [3:0] MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_1_or_ssc;
  reg [4:0] operator_ac_float_cctor_m_34_lpi_1_dfm_10_6;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_8_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_6_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0;
  reg MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_5;
  reg MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_4;
  reg MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5;
  reg MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_8_ssc;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_9_ssc;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_10_ssc;
  wire or_973_cse;
  wire or_974_cse;
  wire or_985_cse;
  wire or_986_cse;
  wire or_993_cse;
  wire or_994_cse;
  wire or_983_cse;
  wire or_984_cse;
  wire or_991_cse;
  wire or_981_cse;
  wire or_982_cse;
  wire or_989_cse;
  wire or_979_cse;
  wire or_980_cse;
  wire or_977_cse;
  wire or_978_cse;
  wire or_992_cse;
  wire or_975_cse;
  wire or_976_cse;
  wire or_990_cse;
  wire or_987_cse;
  wire or_988_cse;
  wire mux_8_cse;
  wire mux_80_cse;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4;
  wire and_1482_m1c;
  wire and_1486_m1c;
  wire and_1492_m1c;
  wire [4:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  wire [4:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_1_ssc;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0;
  wire [4:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  wire [4:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [4:0] MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  wire [4:0] MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  wire [4:0] MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  wire [4:0] MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb;
  wire [4:0] MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb;
  wire [4:0] MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb;
  wire [4:0] MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb;
  wire [4:0] MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb;
  wire [4:0] MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb;
  wire [4:0] MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb;
  wire [4:0] MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb;
  wire [4:0] MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb;
  wire [4:0] MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb;
  wire [4:0] MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb;
  wire [4:0] MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_10_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_9_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_11_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_13_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_14_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_2_ssc;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse;
  wire and_1587_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_8_cse;
  reg [4:0] delay_lane_imag_e_11_sva;
  reg [4:0] delay_lane_imag_e_14_sva;
  reg [4:0] delay_lane_real_e_2_sva;
  reg [4:0] delay_lane_imag_e_7_sva;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1;
  wire or_dcpl_526;
  wire or_dcpl_527;
  wire or_dcpl_528;
  wire or_dcpl_529;
  wire or_dcpl_530;
  wire or_dcpl_531;
  wire or_dcpl_532;
  wire or_dcpl_533;
  wire or_dcpl_534;
  wire or_dcpl_535;
  wire or_dcpl_536;
  wire or_dcpl_537;
  wire or_dcpl_538;
  wire or_dcpl_539;
  wire or_dcpl_540;
  wire or_dcpl_541;
  wire or_dcpl_543;
  wire or_dcpl_544;
  wire or_dcpl_546;
  wire or_dcpl_548;
  wire or_dcpl_550;
  wire or_dcpl_551;
  wire or_dcpl_552;
  wire or_dcpl_554;
  wire or_dcpl_555;
  wire or_dcpl_558;
  wire or_dcpl_577;
  wire or_dcpl_578;
  wire [4:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [4:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [4:0] MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [4:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire and_1240_ssc;
  wire or_573_ssc;
  wire [4:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [4:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt;
  wire and_1282_ssc;
  wire or_582_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_2_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_3_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_4_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_5_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_6_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_7_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_1_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_2_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_6_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_7_cse;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c6;
  reg [4:0] delay_lane_real_e_10_sva;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  reg [4:0] delay_lane_real_e_11_sva;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2;
  reg [4:0] delay_lane_imag_e_13_sva;
  reg [4:0] delay_lane_real_e_13_sva;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  reg [4:0] delay_lane_imag_e_9_sva;
  reg [4:0] delay_lane_imag_e_10_sva;
  wire [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c5;
  wire [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_3_0;
  wire nor_562_m1c;
  wire nor_561_m1c;
  wire nor_560_m1c;
  wire nor_559_m1c;
  wire nor_558_m1c;
  wire nor_557_m1c;
  wire nor_556_m1c;
  wire nor_555_m1c;
  wire nor_554_m1c;
  wire nor_553_m1c;
  wire nor_552_m1c;
  wire nor_551_m1c;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_ssc;
  wire or_1011_tmp;
  wire or_1065_tmp;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c6;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_4;
  wire [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_3_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_4;
  wire [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_3_0;
  wire [5:0] MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [5:0] MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [6:0] nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [5:0] MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [5:0] MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm;
  wire [6:0] nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm;
  wire [5:0] MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_54_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_57_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_60_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_63_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_66_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_69_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_72_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_35_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_38_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_41_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_44_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_47_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_50_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_3;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_53_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_itm;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_itm;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_3_itm;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_5_itm;
  wire and_1488_itm;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_7_itm;
  wire and_1494_itm;
  wire and_1496_itm;
  wire and_1499_itm;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_itm;
  wire and_1504_itm;
  wire and_1507_itm;
  wire and_1510_itm;
  wire and_1513_itm;
  wire and_1516_itm;
  wire and_1519_itm;
  wire and_1522_itm;
  wire and_1525_itm;
  wire and_1528_itm;
  wire and_1531_itm;
  wire and_1534_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm;
  wire [6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire and_269_itm;
  wire and_272_itm;
  wire and_275_itm;
  wire and_278_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire and_568_itm;
  wire and_571_itm;
  wire and_574_itm;
  wire and_577_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire and_618_itm;
  wire and_621_itm;
  wire and_624_itm;
  wire and_627_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire and_705_itm;
  wire and_708_itm;
  wire and_711_itm;
  wire and_714_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [12:0] MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire and_784_itm;
  wire and_787_itm;
  wire and_790_itm;
  wire and_793_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire and_870_itm;
  wire and_873_itm;
  wire and_876_itm;
  wire and_879_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire and_1318_itm;
  wire and_1321_itm;
  wire and_1324_itm;
  wire and_1327_itm;
  wire [6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [11:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [11:0] MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [12:0] nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [12:0] MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire and_631_itm;
  wire and_634_itm;
  wire and_636_itm;
  wire and_640_itm;
  wire and_642_itm;
  wire nor_270_itm;
  wire and_647_itm;
  wire nor_286_itm;
  wire and_652_itm;
  wire and_655_itm;
  wire and_660_itm;
  wire and_663_itm;
  wire and_666_itm;
  wire and_670_itm;
  wire and_674_itm;
  wire and_677_itm;
  wire and_680_itm;
  wire and_684_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [12:0] MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm;
  wire [12:0] MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_itm;
  wire [12:0] MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_itm;
  wire [5:0] MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm;
  wire [6:0] nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm;
  wire mux_119_itm;
  wire mux_123_itm;
  wire mux_184_itm;
  wire [5:0] z_out;
  wire [6:0] nl_z_out;
  wire [5:0] z_out_1;
  wire [6:0] nl_z_out_1;
  wire [5:0] z_out_2;
  wire [6:0] nl_z_out_2;
  wire [5:0] z_out_3;
  wire [6:0] nl_z_out_3;
  wire and_dcpl_1740;
  wire [6:0] z_out_4;
  wire and_dcpl_1752;
  wire [6:0] z_out_5;
  wire and_dcpl_1779;
  wire and_dcpl_1780;
  wire and_dcpl_1788;
  wire [5:0] z_out_6;
  wire [6:0] z_out_7;
  wire [6:0] z_out_8;
  wire [6:0] z_out_9;
  wire [6:0] z_out_10;
  wire and_dcpl_1857;
  wire and_dcpl_1860;
  wire [6:0] z_out_11;
  wire and_dcpl_1872;
  wire and_dcpl_1875;
  wire [6:0] z_out_12;
  wire and_dcpl_1885;
  wire and_dcpl_1892;
  wire [6:0] z_out_14;
  wire [6:0] z_out_15;
  wire and_dcpl_1939;
  wire and_dcpl_1942;
  wire [6:0] z_out_16;
  wire and_dcpl_1952;
  wire and_dcpl_1962;
  wire [6:0] z_out_18;
  wire [6:0] z_out_19;
  wire [6:0] z_out_20;
  wire and_dcpl_1995;
  wire and_dcpl_1998;
  wire [6:0] z_out_21;
  wire [6:0] z_out_22;
  wire [6:0] z_out_23;
  wire and_dcpl_2029;
  wire [6:0] z_out_25;
  wire [6:0] z_out_26;
  wire [6:0] z_out_27;
  wire [5:0] z_out_28;
  wire [6:0] nl_z_out_28;
  wire [5:0] z_out_29;
  wire [6:0] nl_z_out_29;
  wire [5:0] z_out_30;
  wire [6:0] nl_z_out_30;
  wire [4:0] z_out_31;
  wire [11:0] z_out_33;
  wire [11:0] z_out_34;
  wire [11:0] z_out_35;
  wire [11:0] z_out_36;
  wire [11:0] z_out_37;
  wire [11:0] z_out_38;
  wire [12:0] nl_z_out_38;
  wire [11:0] z_out_39;
  wire [12:0] nl_z_out_39;
  wire [11:0] z_out_40;
  wire [12:0] nl_z_out_40;
  wire [11:0] z_out_41;
  wire [12:0] nl_z_out_41;
  wire [12:0] z_out_42;
  wire [12:0] z_out_43;
  wire [12:0] z_out_44;
  wire [12:0] z_out_45;
  wire [12:0] z_out_46;
  wire [12:0] z_out_47;
  wire [12:0] z_out_48;
  wire [12:0] z_out_49;
  wire [12:0] z_out_50;
  wire [12:0] z_out_51;
  wire [12:0] z_out_52;
  wire [12:0] z_out_53;
  wire [12:0] z_out_54;
  wire [12:0] z_out_55;
  wire [12:0] z_out_56;
  wire [12:0] z_out_57;
  wire [12:0] z_out_58;
  wire [12:0] z_out_59;
  wire [12:0] z_out_60;
  wire [12:0] z_out_61;
  wire [12:0] z_out_62;
  wire [12:0] z_out_63;
  wire [12:0] z_out_64;
  wire [12:0] z_out_65;
  wire [12:0] z_out_66;
  wire [12:0] z_out_67;
  wire [11:0] z_out_68;
  wire and_dcpl_2475;
  wire [11:0] z_out_69;
  wire [11:0] z_out_70;
  reg [4:0] delay_lane_real_e_7_sva;
  reg [4:0] delay_lane_real_e_8_sva;
  reg [4:0] delay_lane_real_e_6_sva;
  reg [4:0] delay_lane_real_e_9_sva;
  reg [4:0] delay_lane_real_e_5_sva;
  reg [4:0] delay_lane_real_e_4_sva;
  reg [4:0] delay_lane_real_e_3_sva;
  reg [4:0] delay_lane_real_e_12_sva;
  reg [4:0] delay_lane_real_e_1_sva;
  reg [4:0] delay_lane_real_e_14_sva;
  reg [4:0] delay_lane_real_e_0_sva;
  reg [4:0] delay_lane_imag_e_8_sva;
  reg [4:0] delay_lane_imag_e_6_sva;
  reg [4:0] delay_lane_imag_e_5_sva;
  reg [4:0] delay_lane_imag_e_4_sva;
  reg [4:0] delay_lane_imag_e_3_sva;
  reg [4:0] delay_lane_imag_e_12_sva;
  reg [4:0] delay_lane_imag_e_2_sva;
  reg [4:0] delay_lane_imag_e_1_sva;
  reg [4:0] delay_lane_imag_e_0_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva;
  reg [4:0] operator_ac_float_cctor_e_31_lpi_1_dfm;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva;
  reg [4:0] operator_ac_float_cctor_e_61_lpi_1_dfm;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva;
  reg [4:0] operator_ac_float_cctor_e_62_lpi_1_dfm;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva;
  reg [4:0] operator_ac_float_cctor_e_33_lpi_1_dfm;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva;
  reg [4:0] operator_ac_float_cctor_e_63_lpi_1_dfm;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva;
  reg [4:0] operator_ac_float_cctor_e_34_lpi_1_dfm;
  reg [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  reg [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva;
  reg MAC_1_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_1_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_1_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_1_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_2_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_2_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_2_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_2_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_3_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_3_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_3_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_3_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_4_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_4_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_4_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_4_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_5_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_6_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_6_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_6_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_7_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_7_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_7_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_7_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_8_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_8_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_8_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_8_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_9_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_9_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_9_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_9_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_13_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_13_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_13_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_13_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_14_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_14_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_14_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_14_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_15_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_15_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_15_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_15_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  reg MAC_16_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  reg MAC_16_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  reg MAC_16_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  reg MAC_16_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  wire return_imag_e_rsci_idat_mx0c1;
  wire return_real_e_rsci_idat_mx0c1;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1;
  wire [5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [6:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1;
  wire [5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire [6:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_mx0c2;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_mx0w2;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c9;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c10;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c11;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c12;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c13;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c14;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c15;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c16;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c17;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c18;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c19;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c20;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c21;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c22;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c23;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c7;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c8;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c4;
  wire my_complex_float_t_cctor_imag_operator_return_4_sva_mx0w1;
  wire my_complex_float_t_cctor_real_operator_return_9_sva_mx0w1;
  wire my_complex_float_t_cctor_imag_operator_return_3_sva_mx0w3;
  wire my_complex_float_t_cctor_imag_operator_return_13_sva_mx0w2;
  wire my_complex_float_t_cctor_imag_operator_return_14_sva_mx0w2;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_itm_mx0w7;
  wire my_complex_float_t_cctor_imag_operator_return_sva_mx0w6;
  wire my_complex_float_t_cctor_real_operator_return_10_sva_mx0w6;
  wire my_complex_float_t_cctor_real_operator_return_11_sva_mx0w5;
  wire my_complex_float_t_cctor_real_operator_return_12_sva_mx0w5;
  wire my_complex_float_t_cctor_real_operator_return_4_sva_mx0w5;
  wire operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c4;
  wire operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c4;
  wire operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c4;
  wire operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c4;
  wire operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c3;
  wire operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c1;
  wire operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c2;
  wire operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c3;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1;
  wire [4:0] operator_ac_float_cctor_e_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_1_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1;
  wire [4:0] operator_ac_float_cctor_e_13_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_28_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1;
  wire [4:0] operator_ac_float_cctor_e_12_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_27_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1;
  wire [4:0] operator_ac_float_cctor_e_11_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_26_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1;
  wire [4:0] operator_ac_float_cctor_e_10_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_25_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_9_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_24_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1;
  wire [4:0] operator_ac_float_cctor_e_8_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_23_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1;
  wire [4:0] operator_ac_float_cctor_e_7_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_22_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1;
  wire [4:0] operator_ac_float_cctor_e_21_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0;
  wire [1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
  wire [2:0] nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
  wire [1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
  wire [2:0] nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
  wire [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_16_sva_1;
  wire [4:0] operator_ac_float_cctor_e_15_lpi_1_dfm_mx0;
  wire [4:0] operator_ac_float_cctor_e_30_lpi_1_dfm_mx0;
  wire [11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1;
  wire [12:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1;
  wire [12:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_mx0w0;
  wire [3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0;
  wire [3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0;
  reg MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_4;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_4;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_70;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_105;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_71;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_106;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_72;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_107;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_73;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_108;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_74;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_109;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_75;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_110;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_76;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_111;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_77;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_112;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_78;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_113;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_79;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_114;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_80;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_115;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_81;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_116;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_82;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_117;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_83;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_118;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_84;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_119;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_85;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_120;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_86;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_121;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_87;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_122;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_88;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_123;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_89;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_124;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_90;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_125;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_91;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_126;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_92;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_127;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_93;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_128;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_94;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_129;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_95;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_130;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_96;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_131;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_97;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_132;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_98;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_133;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_99;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_134;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_100;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_135;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_101;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_136;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_102;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_137;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_103;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_138;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_104;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_139;
  wire [4:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_conc_32_itm_4_0;
  wire [4:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_conc_29_itm_4_0;
  wire [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0;
  wire [6:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0;
  wire [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0;
  wire [6:0] nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0;
  wire [5:0] ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0;
  wire [6:0] nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0;
  wire [5:0] ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0;
  wire [6:0] nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2;
  reg [1:0] operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0;
  reg [3:0] operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1;
  reg [4:0] operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0;
  reg [1:0] operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1;
  reg [3:0] operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0;
  reg [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_1_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_2_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_26_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_27_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_28_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_29_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_30_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_31_ssc;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0;
  reg [5:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_2_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_3_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_4_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_5_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_6_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_7_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_2_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_3_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_4_ssc;
  reg [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_5_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_ssc;
  reg [3:0] operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_1_ssc;
  reg [3:0] operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_6_ssc;
  reg [3:0] operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_7_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_54_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_55_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_28_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_44_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_5_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_11_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_62_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_63_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_50_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_51_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_26_ssc;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_42_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_58_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_59_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_62_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_63_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_58_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_59_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_30_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_31_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_26_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_27_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_22_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_23_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_22_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_23_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_18_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_19_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_18_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_19_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_10_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_11_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_6_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_7_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_2_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_3_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_46_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_47_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_42_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_43_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_39_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_39_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_38_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_39_ssc;
  wire and_1785_m1c;
  wire [4:0] operator_r_m_6_lpi_1_dfm_mx0w5_10_6;
  wire [4:0] operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_10_6;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_10_6;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_15_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_10_6;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_14_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_10_6;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_13_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_10_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_10_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_10_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_8_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_8_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_7_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_6_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_6_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_5_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_5_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_4_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_4_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_3_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_2_lpi_1_dfm_1_5_0;
  wire [4:0] operator_i_m_8_lpi_1_dfm_mx0w10_10_6;
  wire [4:0] operator_i_m_7_lpi_1_dfm_mx0w3_10_6;
  wire [4:0] operator_i_m_6_lpi_1_dfm_mx0w4_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_2_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6;
  wire [4:0] operator_r_m_3_lpi_1_dfm_mx0w6_10_6;
  wire [4:0] operator_r_m_2_lpi_1_dfm_mx0w6_10_6;
  wire [4:0] operator_i_m_9_lpi_1_dfm_mx0w10_10_6;
  wire [4:0] operator_r_m_lpi_1_dfm_mx0w6_10_6;
  wire and_594_ssc;
  wire and_597_ssc;
  wire and_606_ssc;
  wire and_609_ssc;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0;
  wire [4:0] operator_r_m_15_lpi_1_dfm_mx0w4_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_1_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_5_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_4_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1_4_0;
  wire [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_4_0;
  wire [4:0] operator_i_m_1_lpi_1_dfm_mx0w3_10_6;
  wire [5:0] operator_i_m_1_lpi_1_dfm_mx0w3_5_0;
  wire [4:0] operator_ac_float_cctor_m_1_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_35_lpi_1_dfm_1_10_6;
  wire [5:0] operator_ac_float_cctor_m_35_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_28_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_27_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_41_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_26_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_40_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_25_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_24_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_23_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_22_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_21_lpi_1_dfm_1_10_6;
  wire [5:0] operator_ac_float_cctor_m_21_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_47_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_46_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_45_lpi_1_dfm_1_10_6;
  wire [5:0] operator_ac_float_cctor_m_45_lpi_1_dfm_1_5_0;
  wire [4:0] operator_ac_float_cctor_m_60_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_30_lpi_1_dfm_1_10_6;
  wire [5:0] operator_ac_float_cctor_m_30_lpi_1_dfm_1_5_0;
  wire [5:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt;
  wire [6:0] nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt;
  wire [5:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt;
  wire [6:0] nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt;
  wire [5:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt;
  wire [6:0] nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt;
  wire [5:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt;
  wire [6:0] nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt;
  wire [5:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt;
  wire [6:0] nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt;
  wire [6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt;
  wire [7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire [7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire [6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt;
  wire [6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire [7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  wire [4:0] operator_r_m_4_lpi_1_dfm_mx0w5_10_6;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  wire [3:0] operator_r_m_14_lpi_1_dfm_mx0w5_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_9_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_7_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_6_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_5_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_3_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_2_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_2_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_1_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6;
  wire and_537_ssc;
  wire and_540_ssc;
  wire and_543_ssc;
  wire and_546_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_ssc;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6;
  reg [4:0] operator_ac_float_cctor_m_63_lpi_1_dfm_10_6;
  reg [4:0] operator_ac_float_cctor_m_64_lpi_1_dfm_10_6;
  reg [4:0] operator_ac_float_cctor_m_65_lpi_1_dfm_10_6;
  wire [4:0] operator_r_m_1_lpi_1_dfm_mx0w4_10_6;
  wire [5:0] operator_r_m_1_lpi_1_dfm_mx0w4_5_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_30_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_31_ssc;
  wire [4:0] operator_ac_float_cctor_m_43_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_26_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_27_ssc;
  wire [4:0] operator_ac_float_cctor_m_42_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_14_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_15_ssc;
  wire [3:0] operator_ac_float_cctor_m_54_lpi_1_dfm_1_3_0;
  wire nor_501_cse;
  wire nor_578_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse;
  wire and_969_rgt;
  wire or_487_rgt;
  wire and_1331_rgt;
  wire or_590_rgt;
  wire or_736_rgt;
  wire and_1462_rgt;
  wire and_1465_rgt;
  wire and_1466_rgt;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1;
  reg [4:0] operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0;
  reg [1:0] operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1;
  reg [4:0] operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0;
  reg [1:0] operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1;
  reg [4:0] operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0;
  reg [1:0] operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_8_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_17_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_10_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_11_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_10_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_11_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_6_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_7_ssc;
  wire nor_474_tmp;
  wire nor_495_tmp;
  wire nor_493_tmp;
  wire nor_489_tmp;
  wire nor_487_tmp;
  wire nor_485_tmp;
  wire nor_519_tmp;
  wire nor_491_tmp;
  wire nor_476_tmp;
  wire [4:0] operator_r_m_9_lpi_1_dfm_mx0w6_10_6;
  wire [4:0] operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_8_ssc;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_4_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_1_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_ssc;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_3_0;
  wire and_462_ssc;
  wire and_465_ssc;
  wire and_468_ssc;
  wire and_471_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_7_ssc;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6;
  wire [4:0] operator_ac_float_cctor_m_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_38_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_53_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6;
  wire [6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire [7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt;
  wire [6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire [7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0;
  wire [1:0] operator_r_m_3_lpi_1_dfm_mx0w6_5_4;
  wire [3:0] operator_r_m_3_lpi_1_dfm_mx0w6_3_0;
  wire [1:0] operator_r_m_2_lpi_1_dfm_mx0w6_5_4;
  wire [3:0] operator_r_m_2_lpi_1_dfm_mx0w6_3_0;
  wire [1:0] operator_r_m_lpi_1_dfm_mx0w6_5_4;
  wire [3:0] operator_r_m_lpi_1_dfm_mx0w6_3_0;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4;
  wire [1:0] operator_r_m_15_lpi_1_dfm_mx0w4_5_4;
  wire [3:0] operator_r_m_15_lpi_1_dfm_mx0w4_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_41_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_41_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_40_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_40_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_23_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_23_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_22_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_22_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_47_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_47_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_46_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_46_lpi_1_dfm_1_3_0;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_6_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_13_ssc;
  wire [4:0] operator_r_m_7_lpi_1_dfm_mx0w4_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_6_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_5_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6;
  wire and_506_ssc;
  wire and_509_ssc;
  wire and_512_ssc;
  wire and_515_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_8_ssc;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_ssc;
  wire [4:0] operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6;
  wire [11:0] MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire [12:0] nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_6_ssc;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_ssc;
  wire [3:0] operator_ac_float_cctor_m_20_lpi_1_dfm_1_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_6_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_7_ssc;
  wire [4:0] operator_ac_float_cctor_m_52_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_2_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_3_ssc;
  wire [4:0] operator_ac_float_cctor_m_36_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_2_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_3_ssc;
  wire [4:0] operator_ac_float_cctor_m_51_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_ssc;
  wire [3:0] operator_ac_float_cctor_m_6_lpi_1_dfm_1_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_ssc;
  wire [4:0] operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6;
  wire [1:0] operator_r_m_4_lpi_1_dfm_mx0w5_5_4;
  wire [3:0] operator_r_m_4_lpi_1_dfm_mx0w5_3_0;
  wire [4:0] operator_r_m_14_lpi_1_dfm_mx0w5_10_6;
  wire [1:0] operator_r_m_14_lpi_1_dfm_mx0w5_5_4;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_43_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_43_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_42_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_42_lpi_1_dfm_1_3_0;
  wire [4:0] operator_ac_float_cctor_m_54_lpi_1_dfm_1_10_6;
  wire [1:0] operator_ac_float_cctor_m_54_lpi_1_dfm_1_5_4;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0;
  wire and_1893_cse;
  wire and_2125_cse;
  wire and_2241_cse;
  wire and_2326_cse;
  wire and_2317_cse;
  wire and_2438_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_71_cse;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_7_ssc;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_15_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_30_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_31_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_26_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_27_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_6_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_7_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_ssc;
  wire [3:0] operator_r_m_8_lpi_1_dfm_mx0w6_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_4_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_3_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6;
  wire and_581_ssc;
  wire and_584_ssc;
  wire and_587_ssc;
  wire and_590_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_10_ssc;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6;
  wire [4:0] operator_ac_float_cctor_m_58_lpi_1_dfm_1_10_6;
  wire [4:0] operator_ac_float_cctor_m_57_lpi_1_dfm_1_10_6;
  wire [3:0] operator_ac_float_cctor_m_37_lpi_1_dfm_1_3_0;
  wire [3:0] operator_ac_float_cctor_m_17_lpi_1_dfm_1_3_0;
  wire [6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire [7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6;
  wire [6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire [7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_5_4;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_5_4;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_12_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_12_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_11_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_11_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_53_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_53_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_8_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_8_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_7_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_7_lpi_1_dfm_1_3_0;
  reg [4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4;
  wire [1:0] operator_ac_float_cctor_m_52_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_52_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_51_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_51_lpi_1_dfm_1_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_ssc;
  wire [4:0] operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_10_6;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_7_ssc;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_22_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_23_ssc;
  wire [4:0] operator_ac_float_cctor_m_56_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_18_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_19_ssc;
  wire [4:0] operator_ac_float_cctor_m_55_lpi_1_dfm_1_10_6;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_14_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_15_ssc;
  wire [4:0] operator_ac_float_cctor_m_39_lpi_1_dfm_1_10_6;
  wire [1:0] operator_r_m_7_lpi_1_dfm_mx0w4_5_4;
  wire [3:0] operator_r_m_7_lpi_1_dfm_mx0w4_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_3_0;
  wire [4:0] operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6;
  wire [1:0] operator_ac_float_cctor_m_20_lpi_1_dfm_1_5_4;
  wire [1:0] operator_ac_float_cctor_m_36_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_36_lpi_1_dfm_1_3_0;
  wire [4:0] operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6;
  wire [1:0] operator_ac_float_cctor_m_6_lpi_1_dfm_1_5_4;
  wire [1:0] operator_ac_float_cctor_m_16_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_16_lpi_1_dfm_1_3_0;
  wire [4:0] operator_r_m_8_lpi_1_dfm_mx0w6_10_6;
  wire [1:0] operator_r_m_8_lpi_1_dfm_mx0w6_5_4;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_3_0;
  wire [4:0] operator_ac_float_cctor_m_37_lpi_1_dfm_1_10_6;
  wire [1:0] operator_ac_float_cctor_m_37_lpi_1_dfm_1_5_4;
  wire [4:0] operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6;
  wire [1:0] operator_ac_float_cctor_m_17_lpi_1_dfm_1_5_4;
  wire and_1886_cse;
  wire and_1888_cse;
  wire and_1899_cse;
  wire and_1909_cse;
  wire and_1883_cse;
  wire and_1925_cse;
  wire and_2261_cse;
  wire and_2264_cse;
  wire reg_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_1_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_5_cse;
  wire [6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_seb;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6;
  wire [6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire [7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_58_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_58_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_57_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_57_lpi_1_dfm_1_3_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4;
  wire [1:0] operator_ac_float_cctor_m_56_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_56_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_55_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_55_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_ac_float_cctor_m_39_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_39_lpi_1_dfm_1_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_90_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_1_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_cse;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_10_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_10_lpi_1_dfm_1_3_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_12_cse;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_6_cse;
  wire not_tmp_1312;
  wire not_tmp_1322;
  wire nor_cse;
  wire or_1078_cse;
  wire and_2663_cse;
  wire nor_536_cse;
  wire nor_534_cse;
  wire nor_774_cse;
  wire mux_561_cse;
  wire nor_794_cse;
  wire nor_796_cse;
  wire mux_536_cse;
  wire [6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_itm;
  wire [5:0] and_1787_itm;
  wire [5:0] MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [6:0] nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [5:0] MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [6:0] nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [5:0] MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm;
  wire [6:0] nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm;
  wire [5:0] MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [6:0] nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm;
  wire [5:0] MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [6:0] nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm;
  wire [5:0] MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [6:0] nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm;
  wire [6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_itm;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_itm;
  wire [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_itm;
  wire [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_itm;
  wire [4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_itm;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  wire MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  wire MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6;
  wire MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1;
  wire MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_4_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_5_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_7_ssc;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_8_ssc;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_6_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_7_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0;
  reg [5:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_8_ssc;
  reg ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_9_ssc;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1;
  reg [1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0;
  reg [3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1;
  wire or_805_ssc;
  wire or_806_ssc;
  wire or_865_ssc;
  wire [4:0] MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [4:0] MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire [5:0] nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_21_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_11_ssc;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_8_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_1_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_3_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_ssc;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_13_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_31_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_33_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_35_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_5_ssc;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0;
  wire operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_4;
  wire [3:0] operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_3_0;
  wire operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_4;
  wire [3:0] operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_3_0;
  wire operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_4;
  wire [3:0] operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_3_0;
  wire [1:0] operator_r_m_6_lpi_1_dfm_mx0w5_5_4;
  wire [3:0] operator_r_m_6_lpi_1_dfm_mx0w5_3_0;
  wire [1:0] operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_5_4;
  wire [3:0] operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_3_0;
  wire [1:0] operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_i_m_8_lpi_1_dfm_mx0w10_5_4;
  wire [3:0] operator_i_m_8_lpi_1_dfm_mx0w10_3_0;
  wire [1:0] operator_i_m_7_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_i_m_7_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_i_m_6_lpi_1_dfm_mx0w4_5_4;
  wire [3:0] operator_i_m_6_lpi_1_dfm_mx0w4_3_0;
  wire [1:0] operator_i_m_9_lpi_1_dfm_mx0w10_5_4;
  wire [3:0] operator_i_m_9_lpi_1_dfm_mx0w10_3_0;
  wire [1:0] operator_ac_float_cctor_m_1_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_1_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_28_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_28_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_27_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_27_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_26_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_26_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_25_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_25_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_24_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_24_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_60_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_60_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_15_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_15_lpi_1_dfm_1_3_0;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_31_ssc;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_32_ssc;
  reg operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0;
  reg [1:0] operator_ac_float_cctor_m_63_lpi_1_dfm_5_4;
  reg [3:0] operator_ac_float_cctor_m_63_lpi_1_dfm_3_0;
  reg [1:0] operator_ac_float_cctor_m_64_lpi_1_dfm_5_4;
  reg [3:0] operator_ac_float_cctor_m_64_lpi_1_dfm_3_0;
  reg [1:0] operator_ac_float_cctor_m_65_lpi_1_dfm_5_4;
  reg [3:0] operator_ac_float_cctor_m_65_lpi_1_dfm_3_0;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_33_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_35_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_38_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_41_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_44_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_46_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_48_cse;
  wire [1:0] operator_r_m_9_lpi_1_dfm_mx0w6_5_4;
  wire [3:0] operator_r_m_9_lpi_1_dfm_mx0w6_3_0;
  wire [1:0] operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_5_4;
  wire [3:0] operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_3_0;
  wire [1:0] operator_ac_float_cctor_m_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_13_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_13_lpi_1_dfm_1_3_0;
  wire [1:0] operator_ac_float_cctor_m_38_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_38_lpi_1_dfm_1_3_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0;
  wire [1:0] operator_ac_float_cctor_m_9_lpi_1_dfm_1_5_4;
  wire [3:0] operator_ac_float_cctor_m_9_lpi_1_dfm_1_3_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc;
  wire z_out_32_4;
  wire [3:0] z_out_32_3_0;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_38_tmp;

  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_1_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_2_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_3_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_1_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_2_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_3_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_1_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_2_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_3_nl;
  wire MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl;
  wire MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl;
  wire MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_4_nl;
  wire MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_5_nl;
  wire MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_6_nl;
  wire MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_7_nl;
  wire MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_4_nl;
  wire MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_5_nl;
  wire MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_6_nl;
  wire MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_7_nl;
  wire MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_4_nl;
  wire MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_5_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_2_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_13_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl;
  wire[3:0] mux1h_12_nl;
  wire and_1233_nl;
  wire and_1236_nl;
  wire and_1239_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_24_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_25_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_26_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_27_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_28_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_29_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_30_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_31_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_32_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_33_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_34_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_35_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_36_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_37_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_38_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_39_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_40_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_41_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_42_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_43_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_44_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_45_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_46_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_47_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_48_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_49_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_50_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_51_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_52_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_53_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_54_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_55_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_56_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_57_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_58_nl;
  wire not_1835_nl;
  wire and_1033_nl;
  wire and_1036_nl;
  wire and_1039_nl;
  wire and_951_nl;
  wire and_954_nl;
  wire and_957_nl;
  wire mux_352_nl;
  wire mux_351_nl;
  wire mux_350_nl;
  wire and_972_nl;
  wire and_975_nl;
  wire and_978_nl;
  wire and_1043_nl;
  wire and_1046_nl;
  wire and_1049_nl;
  wire and_1150_nl;
  wire and_1153_nl;
  wire and_1156_nl;
  wire and_1198_nl;
  wire and_1201_nl;
  wire and_1204_nl;
  wire and_1243_nl;
  wire and_1246_nl;
  wire and_1249_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_16_nl;
  wire or_4_nl;
  wire[5:0] MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire mux_110_nl;
  wire mux_109_nl;
  wire mux_108_nl;
  wire[5:0] MAC_10_r_ac_float_2_else_and_nl;
  wire[1:0] MAC_11_r_ac_float_2_else_and_nl;
  wire[3:0] MAC_11_r_ac_float_2_else_and_1_nl;
  wire[5:0] MAC_12_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_13_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_14_r_ac_float_2_else_and_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_17_nl;
  wire mux_537_nl;
  wire mux_535_nl;
  wire or_1077_nl;
  wire[5:0] and_1827_nl;
  wire[5:0] mux1h_nl;
  wire[5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire and_1832_nl;
  wire and_1833_nl;
  wire not_1834_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_18_nl;
  wire[5:0] and_1820_nl;
  wire[5:0] mux1h_1_nl;
  wire[5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire and_1825_nl;
  wire and_1826_nl;
  wire not_1833_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_19_nl;
  wire[5:0] and_1813_nl;
  wire[5:0] mux1h_2_nl;
  wire[5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire and_1818_nl;
  wire and_1819_nl;
  wire not_1832_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_16_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_17_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_18_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_41_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_19_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_45_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_20_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_49_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_21_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_53_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_22_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_57_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_16_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_61_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_17_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_37_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_18_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_19_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_20_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_21_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_22_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_20_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_21_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_22_nl;
  wire[7:0] acc_17_nl;
  wire[8:0] nl_acc_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_4_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl;
  wire[7:0] acc_13_nl;
  wire[8:0] nl_acc_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_3_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_30_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_15_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_28_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_14_nl;
  wire mux_509_nl;
  wire mux_508_nl;
  wire mux_507_nl;
  wire mux_506_nl;
  wire mux_505_nl;
  wire nor_502_nl;
  wire nor_504_nl;
  wire and_1630_nl;
  wire mux_504_nl;
  wire mux_503_nl;
  wire nor_505_nl;
  wire nor_506_nl;
  wire mux_502_nl;
  wire nor_507_nl;
  wire nor_508_nl;
  wire mux_501_nl;
  wire mux_500_nl;
  wire mux_499_nl;
  wire nor_509_nl;
  wire nor_510_nl;
  wire mux_498_nl;
  wire nor_511_nl;
  wire nor_512_nl;
  wire mux_497_nl;
  wire mux_496_nl;
  wire nor_513_nl;
  wire nor_514_nl;
  wire mux_495_nl;
  wire nor_515_nl;
  wire nor_516_nl;
  wire mux_486_nl;
  wire mux_485_nl;
  wire or_761_nl;
  wire mux_484_nl;
  wire mux_492_nl;
  wire mux_491_nl;
  wire mux_490_nl;
  wire or_765_nl;
  wire or_764_nl;
  wire mux_494_nl;
  wire mux_493_nl;
  wire nor_498_nl;
  wire nor_499_nl;
  wire nor_500_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_nl;
  wire[7:0] acc_24_nl;
  wire[8:0] nl_acc_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_5_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl;
  wire[5:0] and_1779_nl;
  wire[5:0] mux1h_8_nl;
  wire[5:0] MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire and_1782_nl;
  wire and_1783_nl;
  wire and_1784_nl;
  wire or_nl;
  wire and_2626_nl;
  wire not_1826_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl;
  wire[5:0] and_1771_nl;
  wire[5:0] mux1h_9_nl;
  wire[5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire or_1074_nl;
  wire or_1075_nl;
  wire not_1825_nl;
  wire[5:0] MAC_13_r_ac_float_3_else_and_nl;
  wire[5:0] MAC_14_r_ac_float_3_else_and_nl;
  wire mux_198_nl;
  wire mux_197_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire mux_205_nl;
  wire mux_204_nl;
  wire mux_203_nl;
  wire mux_575_nl;
  wire mux_214_nl;
  wire mux_213_nl;
  wire mux_212_nl;
  wire mux_211_nl;
  wire mux_221_nl;
  wire mux_220_nl;
  wire mux_219_nl;
  wire mux_226_nl;
  wire nor_235_nl;
  wire mux_225_nl;
  wire MAC_9_r_ac_float_1_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_1_else_and_1_nl;
  wire mux_234_nl;
  wire or_378_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_7_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_16_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl;
  wire mux_482_nl;
  wire mux_481_nl;
  wire nand_54_nl;
  wire or_744_nl;
  wire or_742_nl;
  wire mux_480_nl;
  wire or_741_nl;
  wire nor_71_nl;
  wire and_1469_nl;
  wire and_1472_nl;
  wire and_1473_nl;
  wire[4:0] result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl;
  wire[5:0] result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl;
  wire result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl;
  wire[4:0] result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[5:0] result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl;
  wire[4:0] result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl;
  wire[5:0] result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl;
  wire[4:0] result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[5:0] result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl;
  wire[5:0] MAC_13_r_ac_float_4_else_and_nl;
  wire[5:0] MAC_14_r_ac_float_4_else_and_nl;
  wire[5:0] MAC_15_r_ac_float_4_else_and_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl;
  wire mux_270_nl;
  wire and_1610_nl;
  wire nor_265_nl;
  wire mux_271_nl;
  wire nor_266_nl;
  wire mux_272_nl;
  wire nor_267_nl;
  wire nor_268_nl;
  wire mux_273_nl;
  wire nand_44_nl;
  wire or_904_nl;
  wire mux_287_nl;
  wire mux_286_nl;
  wire mux_285_nl;
  wire or_905_nl;
  wire mux_284_nl;
  wire or_906_nl;
  wire or_907_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire or_908_nl;
  wire or_909_nl;
  wire mux_281_nl;
  wire or_910_nl;
  wire or_911_nl;
  wire mux_280_nl;
  wire mux_279_nl;
  wire mux_278_nl;
  wire or_912_nl;
  wire or_913_nl;
  wire mux_277_nl;
  wire or_914_nl;
  wire or_915_nl;
  wire mux_276_nl;
  wire mux_275_nl;
  wire or_916_nl;
  wire or_917_nl;
  wire mux_274_nl;
  wire or_918_nl;
  wire or_919_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_28_nl;
  wire[4:0] MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_7_nl;
  wire[4:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_5_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_3_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_15_nl;
  wire[3:0] nor_566_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_16_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_17_nl;
  wire or_1068_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_11_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_39_nl;
  wire[4:0] MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_nl;
  wire MAC_11_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl;
  wire MAC_16_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire MAC_12_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl;
  wire MAC_13_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl;
  wire MAC_14_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl;
  wire MAC_11_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_1_nl;
  wire MAC_12_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_2_nl;
  wire MAC_13_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_3_nl;
  wire MAC_14_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_4_nl;
  wire MAC_15_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl;
  wire MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl;
  wire or_897_nl;
  wire MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_1_nl;
  wire MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl;
  wire or_899_nl;
  wire MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl;
  wire MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl;
  wire MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_1_nl;
  wire MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_10_nl;
  wire MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_11_nl;
  wire MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_12_nl;
  wire MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_13_nl;
  wire MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_2_nl;
  wire MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_3_nl;
  wire or_898_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_9_nl;
  wire MAC_6_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_4_nl;
  wire MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl;
  wire MAC_7_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_5_nl;
  wire MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl;
  wire MAC_8_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_6_nl;
  wire MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl;
  wire MAC_9_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_15_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_15_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_14_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl;
  wire result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl;
  wire[3:0] mux1h_13_nl;
  wire and_960_nl;
  wire and_963_nl;
  wire and_966_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_3_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_5_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_6_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_9_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_10_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_12_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_16_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_17_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_18_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_19_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_20_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_21_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_22_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_24_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_25_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_26_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_27_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_28_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_29_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_30_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_31_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_32_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_33_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_34_nl;
  wire not_1837_nl;
  wire mux_355_nl;
  wire mux_354_nl;
  wire mux_353_nl;
  wire or_486_nl;
  wire[4:0] MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_38_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_16_nl;
  wire mux_443_nl;
  wire mux_442_nl;
  wire nor_138_nl;
  wire mux_400_nl;
  wire mux_396_nl;
  wire mux_395_nl;
  wire nor_53_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_6_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_8_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_13_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_36_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_82_nl;
  wire mux_449_nl;
  wire mux_448_nl;
  wire mux_447_nl;
  wire or_707_nl;
  wire mux_246_nl;
  wire mux_245_nl;
  wire or_392_nl;
  wire mux_454_nl;
  wire mux_453_nl;
  wire mux_452_nl;
  wire mux_451_nl;
  wire mux_251_nl;
  wire mux_250_nl;
  wire mux_249_nl;
  wire mux_463_nl;
  wire nor_205_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire or_399_nl;
  wire[1:0] MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_4_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_5_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_28_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_29_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_40_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_41_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_24_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_25_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_38_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_20_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_21_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_36_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_16_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_17_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_12_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_13_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_39_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_8_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_9_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_37_nl;
  wire[5:0] MAC_2_r_ac_float_4_else_and_nl;
  wire MAC_3_r_ac_float_4_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_4_else_and_1_nl;
  wire MAC_4_r_ac_float_4_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_4_else_and_1_nl;
  wire MAC_5_r_ac_float_4_else_and_nl;
  wire MAC_5_r_ac_float_4_else_and_1_nl;
  wire[3:0] MAC_5_r_ac_float_4_else_and_2_nl;
  wire MAC_3_r_ac_float_2_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_2_else_and_1_nl;
  wire MAC_4_r_ac_float_2_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_2_else_and_1_nl;
  wire MAC_5_r_ac_float_2_else_and_nl;
  wire MAC_5_r_ac_float_2_else_and_1_nl;
  wire[3:0] MAC_5_r_ac_float_2_else_and_2_nl;
  wire[1:0] MAC_6_r_ac_float_2_else_and_nl;
  wire[3:0] MAC_6_r_ac_float_2_else_and_1_nl;
  wire[1:0] MAC_7_r_ac_float_2_else_and_nl;
  wire[3:0] MAC_7_r_ac_float_2_else_and_1_nl;
  wire[5:0] MAC_8_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_16_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_2_r_ac_float_3_else_and_nl;
  wire MAC_3_r_ac_float_3_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_3_else_and_1_nl;
  wire MAC_4_r_ac_float_3_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_3_else_and_1_nl;
  wire MAC_5_r_ac_float_3_else_and_nl;
  wire MAC_5_r_ac_float_3_else_and_1_nl;
  wire[3:0] MAC_5_r_ac_float_3_else_and_2_nl;
  wire MAC_6_r_ac_float_3_else_and_nl;
  wire MAC_6_r_ac_float_3_else_and_1_nl;
  wire[3:0] MAC_6_r_ac_float_3_else_and_2_nl;
  wire[1:0] MAC_7_r_ac_float_3_else_and_nl;
  wire[3:0] MAC_7_r_ac_float_3_else_and_1_nl;
  wire[5:0] MAC_8_r_ac_float_3_else_and_nl;
  wire[5:0] MAC_6_r_ac_float_4_else_and_nl;
  wire[5:0] MAC_7_r_ac_float_4_else_and_nl;
  wire[5:0] MAC_8_r_ac_float_4_else_and_nl;
  wire MAC_3_r_ac_float_1_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_1_else_and_1_nl;
  wire MAC_4_r_ac_float_1_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_1_else_and_1_nl;
  wire[5:0] MAC_6_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_7_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_8_r_ac_float_1_else_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_55_nl;
  wire[1:0] MAC_5_r_ac_float_1_else_and_nl;
  wire[3:0] MAC_5_r_ac_float_1_else_and_1_nl;
  wire[5:0] MAC_16_r_ac_float_1_else_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_35_nl;
  wire[5:0] MAC_1_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_1_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_1_r_ac_float_3_else_and_nl;
  wire[5:0] MAC_1_r_ac_float_4_else_and_nl;
  wire MAC_2_r_ac_float_1_else_and_nl;
  wire[4:0] MAC_2_r_ac_float_1_else_and_1_nl;
  wire[5:0] MAC_2_r_ac_float_2_else_and_nl;
  wire[5:0] MAC_15_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_15_r_ac_float_2_else_and_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_66_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_86_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_85_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_94_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_68_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_82_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_48_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_17_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_92_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_65_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_83_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_35_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_45_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_34_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_43_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_63_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_47_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_51_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_20_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_27_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_78_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_43_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_47_nl;
  wire[4:0] ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_32_nl;
  wire MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nand_nl;
  wire[3:0] MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nor_nl;
  wire not_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_59_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_55_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_51_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_61_nl;
  wire or_803_nl;
  wire or_804_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_49_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_18_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_57_nl;
  wire ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl;
  wire ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_1_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_35_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_30_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_53_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_53_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_49_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_49_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_45_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_45_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_41_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_41_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_33_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_33_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_33_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_76_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_39_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_95_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_26_nl;
  wire or_812_nl;
  wire or_814_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_50_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_19_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_77_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_40_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_96_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_27_nl;
  wire or_820_nl;
  wire or_822_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_40_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_20_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_93_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_41_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_97_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_32_nl;
  wire or_828_nl;
  wire or_830_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_41_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_21_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_94_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_42_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_33_nl;
  wire or_836_nl;
  wire or_838_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_46_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_29_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_100_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_51_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_103_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_42_nl;
  wire or_844_nl;
  wire or_846_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_51_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_22_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_74_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_56_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_108_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_26_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_36_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_90_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_20_nl;
  wire or_852_nl;
  wire or_854_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_42_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_23_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_43_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_99_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_30_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_73_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_37_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_91_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_23_nl;
  wire or_860_nl;
  wire or_862_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_43_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_24_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_96_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_50_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_101_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_29_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_74_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_38_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_92_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_24_nl;
  wire ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_2_nl;
  wire or_866_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_36_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_31_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_37_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_33_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_44_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_32_nl;
  wire or_887_nl;
  wire or_889_nl;
  wire[6:0] MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[5:0] MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[5:0] MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl;
  wire[7:0] nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl;
  wire[6:0] MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl;
  wire[7:0] nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl;
  wire[5:0] MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire[6:0] nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl;
  wire mux_106_nl;
  wire mux_113_nl;
  wire mux_118_nl;
  wire mux_117_nl;
  wire nand_nl;
  wire mux_116_nl;
  wire mux_115_nl;
  wire mux_114_nl;
  wire mux_122_nl;
  wire or_319_nl;
  wire mux_121_nl;
  wire mux_120_nl;
  wire mux_102_nl;
  wire or_323_nl;
  wire mux_145_nl;
  wire mux_147_nl;
  wire mux_146_nl;
  wire mux_154_nl;
  wire and_245_nl;
  wire mux_161_nl;
  wire or_51_nl;
  wire mux_175_nl;
  wire mux_183_nl;
  wire mux_182_nl;
  wire mux_181_nl;
  wire or_8_nl;
  wire mux_180_nl;
  wire mux_179_nl;
  wire mux_178_nl;
  wire or_57_nl;
  wire nor_177_nl;
  wire or_386_nl;
  wire mux_262_nl;
  wire mux_261_nl;
  wire mux_260_nl;
  wire mux_269_nl;
  wire mux_268_nl;
  wire mux_266_nl;
  wire mux_362_nl;
  wire mux_385_nl;
  wire nor_8_nl;
  wire mux_398_nl;
  wire mux_81_nl;
  wire or_608_nl;
  wire or_760_nl;
  wire mux_488_nl;
  wire or_763_nl;
  wire mux_158_nl;
  wire mux_157_nl;
  wire mux_230_nl;
  wire mux_291_nl;
  wire or_920_nl;
  wire or_921_nl;
  wire mux_292_nl;
  wire nor_295_nl;
  wire nor_296_nl;
  wire mux_306_nl;
  wire mux_305_nl;
  wire mux_304_nl;
  wire or_922_nl;
  wire mux_303_nl;
  wire or_923_nl;
  wire or_924_nl;
  wire mux_302_nl;
  wire mux_301_nl;
  wire or_925_nl;
  wire or_926_nl;
  wire mux_300_nl;
  wire or_927_nl;
  wire or_928_nl;
  wire mux_299_nl;
  wire mux_298_nl;
  wire mux_297_nl;
  wire or_929_nl;
  wire or_930_nl;
  wire mux_296_nl;
  wire or_931_nl;
  wire or_932_nl;
  wire mux_295_nl;
  wire mux_294_nl;
  wire or_933_nl;
  wire or_934_nl;
  wire mux_293_nl;
  wire or_935_nl;
  wire or_936_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire mux_326_nl;
  wire mux_325_nl;
  wire or_937_nl;
  wire or_938_nl;
  wire or_939_nl;
  wire mux_324_nl;
  wire mux_323_nl;
  wire or_940_nl;
  wire or_941_nl;
  wire mux_322_nl;
  wire or_942_nl;
  wire or_943_nl;
  wire mux_321_nl;
  wire mux_320_nl;
  wire mux_319_nl;
  wire or_944_nl;
  wire or_945_nl;
  wire mux_318_nl;
  wire or_946_nl;
  wire or_947_nl;
  wire mux_317_nl;
  wire mux_316_nl;
  wire or_948_nl;
  wire or_949_nl;
  wire mux_315_nl;
  wire or_950_nl;
  wire or_951_nl;
  wire mux_349_nl;
  wire mux_348_nl;
  wire mux_347_nl;
  wire mux_346_nl;
  wire nand_46_nl;
  wire or_952_nl;
  wire or_953_nl;
  wire mux_345_nl;
  wire mux_344_nl;
  wire or_954_nl;
  wire or_955_nl;
  wire mux_343_nl;
  wire or_956_nl;
  wire or_957_nl;
  wire mux_342_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire or_958_nl;
  wire or_959_nl;
  wire mux_339_nl;
  wire or_960_nl;
  wire or_961_nl;
  wire mux_338_nl;
  wire mux_337_nl;
  wire or_962_nl;
  wire or_963_nl;
  wire mux_336_nl;
  wire or_964_nl;
  wire or_965_nl;
  wire mux_360_nl;
  wire nor_389_nl;
  wire mux_359_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire mux_377_nl;
  wire mux_376_nl;
  wire mux_375_nl;
  wire nor_395_nl;
  wire mux_374_nl;
  wire nor_393_nl;
  wire mux_373_nl;
  wire nor_396_nl;
  wire nor_397_nl;
  wire mux_372_nl;
  wire mux_371_nl;
  wire nor_398_nl;
  wire nor_399_nl;
  wire mux_370_nl;
  wire nor_400_nl;
  wire nor_401_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire mux_367_nl;
  wire nor_402_nl;
  wire nor_403_nl;
  wire mux_366_nl;
  wire nor_404_nl;
  wire nor_405_nl;
  wire mux_365_nl;
  wire mux_364_nl;
  wire nor_406_nl;
  wire nor_407_nl;
  wire mux_363_nl;
  wire nor_408_nl;
  wire nor_409_nl;
  wire mux_412_nl;
  wire mux_411_nl;
  wire mux_410_nl;
  wire mux_409_nl;
  wire or_610_nl;
  wire or_609_nl;
  wire or_605_nl;
  wire mux_414_nl;
  wire mux_413_nl;
  wire nor_431_nl;
  wire nor_432_nl;
  wire nor_433_nl;
  wire mux_418_nl;
  wire mux_417_nl;
  wire mux_416_nl;
  wire mux_415_nl;
  wire or_633_nl;
  wire or_632_nl;
  wire or_630_nl;
  wire or_629_nl;
  wire mux_419_nl;
  wire nor_438_nl;
  wire nor_439_nl;
  wire mux_423_nl;
  wire mux_422_nl;
  wire or_652_nl;
  wire mux_421_nl;
  wire mux_420_nl;
  wire or_354_nl;
  wire mux_424_nl;
  wire nor_443_nl;
  wire nor_444_nl;
  wire mux_425_nl;
  wire nor_447_nl;
  wire nor_448_nl;
  wire mux_426_nl;
  wire nor_451_nl;
  wire nor_452_nl;
  wire mux_428_nl;
  wire or_680_nl;
  wire mux_427_nl;
  wire mux_430_nl;
  wire mux_429_nl;
  wire or_687_nl;
  wire or_686_nl;
  wire mux_431_nl;
  wire nor_457_nl;
  wire nor_458_nl;
  wire mux_432_nl;
  wire nor_461_nl;
  wire nor_462_nl;
  wire mux_517_nl;
  wire mux_nl;
  wire or_1030_nl;
  wire mux_518_nl;
  wire nor_567_nl;
  wire nor_568_nl;
  wire mux_519_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_1_nl;
  wire[3:0] nor_574_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_5_nl;
  wire mux_389_nl;
  wire mux_388_nl;
  wire mux_387_nl;
  wire or_572_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire mux_391_nl;
  wire or_581_nl;
  wire mux_528_nl;
  wire mux_527_nl;
  wire mux_526_nl;
  wire mux_533_nl;
  wire[4:0] MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl;
  wire[4:0] MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_39_nl;
  wire[5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire mux_128_nl;
  wire mux_126_nl;
  wire mux_125_nl;
  wire[5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire mux_130_nl;
  wire nor_218_nl;
  wire nor_219_nl;
  wire[5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[5:0] and_1807_nl;
  wire[5:0] mux1h_3_nl;
  wire[5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire and_1811_nl;
  wire and_1812_nl;
  wire not_1831_nl;
  wire[5:0] and_1801_nl;
  wire[5:0] mux1h_4_nl;
  wire[5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire and_1805_nl;
  wire and_1806_nl;
  wire not_1830_nl;
  wire[5:0] and_1795_nl;
  wire[5:0] mux1h_5_nl;
  wire[5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire and_1799_nl;
  wire and_1800_nl;
  wire not_1829_nl;
  wire and_236_nl;
  wire mux_148_nl;
  wire or_337_nl;
  wire mux_551_nl;
  wire[5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_20_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl;
  wire[5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_21_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl;
  wire[5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_22_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl;
  wire[5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_23_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl;
  wire[5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[5:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[5:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[5:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[4:0] MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire mux_150_nl;
  wire[4:0] MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire mux_151_nl;
  wire[4:0] MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl;
  wire[4:0] MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire mux_479_nl;
  wire mux_478_nl;
  wire mux_477_nl;
  wire or_735_nl;
  wire mux_476_nl;
  wire mux_475_nl;
  wire or_733_nl;
  wire mux_474_nl;
  wire mux_473_nl;
  wire mux_472_nl;
  wire or_729_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_33_nl;
  wire[5:0] and_1791_nl;
  wire[5:0] mux1h_6_nl;
  wire[5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire and_1793_nl;
  wire and_1794_nl;
  wire not_1828_nl;
  wire[5:0] mux1h_7_nl;
  wire[5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire and_1789_nl;
  wire and_1790_nl;
  wire not_1827_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl;
  wire mux_553_nl;
  wire mux_552_nl;
  wire or_1097_nl;
  wire or_1094_nl;
  wire or_1093_nl;
  wire or_1091_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl;
  wire mux_555_nl;
  wire or_1109_nl;
  wire mux_554_nl;
  wire or_1108_nl;
  wire or_1105_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_37_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_38_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_22_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_23_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_24_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_25_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_26_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_27_nl;
  wire and_1135_nl;
  wire and_1138_nl;
  wire and_1141_nl;
  wire[5:0] and_1765_nl;
  wire[5:0] mux1h_10_nl;
  wire[5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire[6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl;
  wire or_1076_nl;
  wire and_1770_nl;
  wire not_1824_nl;
  wire[5:0] and_1759_nl;
  wire[5:0] mux1h_11_nl;
  wire[5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire and_1762_nl;
  wire and_1763_nl;
  wire and_1764_nl;
  wire not_1823_nl;
  wire[3:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl;
  wire and_1184_nl;
  wire and_1187_nl;
  wire and_1190_nl;
  wire[5:0] MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire[6:0] nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl;
  wire mux_557_nl;
  wire mux_556_nl;
  wire or_1144_nl;
  wire nor_787_nl;
  wire nor_788_nl;
  wire nor_789_nl;
  wire[5:0] MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire[6:0] nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl;
  wire mux_562_nl;
  wire mux_560_nl;
  wire nor_793_nl;
  wire mux_559_nl;
  wire or_1126_nl;
  wire mux_566_nl;
  wire mux_564_nl;
  wire nor_800_nl;
  wire mux_563_nl;
  wire or_1132_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire mux_288_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire mux_312_nl;
  wire mux_335_nl;
  wire mux_334_nl;
  wire mux_233_nl;
  wire[5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire[6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl;
  wire and_1537_nl;
  wire and_1541_nl;
  wire and_1544_nl;
  wire and_1548_nl;
  wire[5:0] MAC_15_r_ac_float_3_else_and_nl;
  wire[5:0] MAC_16_r_ac_float_3_else_and_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_nl;
  wire[1:0] MAC_10_r_ac_float_4_else_and_nl;
  wire[3:0] MAC_10_r_ac_float_4_else_and_1_nl;
  wire[5:0] MAC_11_r_ac_float_4_else_and_nl;
  wire[5:0] MAC_12_r_ac_float_4_else_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl;
  wire[1:0] MAC_10_r_ac_float_1_else_and_nl;
  wire[3:0] MAC_10_r_ac_float_1_else_and_1_nl;
  wire[5:0] MAC_11_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_12_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_13_r_ac_float_1_else_and_nl;
  wire[5:0] MAC_14_r_ac_float_1_else_and_nl;
  wire mux_569_nl;
  wire mux_568_nl;
  wire mux_567_nl;
  wire and_2677_nl;
  wire and_2678_nl;
  wire nor_751_nl;
  wire nor_807_nl;
  wire nor_808_nl;
  wire nor_809_nl;
  wire and_1285_nl;
  wire and_1288_nl;
  wire and_1291_nl;
  wire and_1334_nl;
  wire and_1337_nl;
  wire and_1340_nl;
  wire and_942_nl;
  wire and_945_nl;
  wire and_948_nl;
  wire mux_460_nl;
  wire mux_459_nl;
  wire mux_458_nl;
  wire nor_470_nl;
  wire mux_256_nl;
  wire mux_255_nl;
  wire mux_254_nl;
  wire mux_252_nl;
  wire[5:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_54_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_nl;
  wire[5:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl;
  wire[1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_71_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_67_nl;
  wire[1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_74_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_68_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_54_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_91_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_80_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_84_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_81_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_49_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_93_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_67_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_75_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_50_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_89_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_76_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_51_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_88_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_77_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_52_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_87_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_78_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_64_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_52_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_104_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_16_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_53_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_90_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_79_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_65_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_55_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_107_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_17_nl;
  wire[1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_73_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_69_nl;
  wire[1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_72_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_70_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_53_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_105_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_18_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_33_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_108_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_64_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_16_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_72_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_48_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_97_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_24_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_65_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_34_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_109_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_17_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_73_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_49_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_25_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_35_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_18_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_67_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_44_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_92_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_19_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_67_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_36_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_111_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_19_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_68_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_45_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_93_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_20_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_68_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_37_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_112_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_20_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_75_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_25_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_64_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_69_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_38_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_113_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_21_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_28_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_104_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_22_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_71_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_29_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_105_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_23_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_72_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_24_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_69_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_46_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_94_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_21_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_47_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_95_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_22_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_71_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_23_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_43_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_99_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_16_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_47_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_73_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_25_nl;
  wire MAC_9_r_ac_float_2_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_2_else_and_1_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_8_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_1_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_1_nl;
  wire[1:0] MAC_10_r_ac_float_3_else_and_nl;
  wire[3:0] MAC_10_r_ac_float_3_else_and_1_nl;
  wire[1:0] MAC_11_r_ac_float_3_else_and_nl;
  wire[3:0] MAC_11_r_ac_float_3_else_and_1_nl;
  wire[5:0] MAC_12_r_ac_float_3_else_and_nl;
  wire[5:0] MAC_16_r_ac_float_4_else_and_nl;
  wire MAC_9_r_ac_float_3_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_3_else_and_1_nl;
  wire MAC_9_r_ac_float_4_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_4_else_and_1_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_38_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_51_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_53_nl;
  wire mux_434_nl;
  wire mux_433_nl;
  wire or_701_nl;
  wire and_1755_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_1_nl;
  wire[3:0] nor_571_nl;
  wire[3:0] nor_572_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_4_nl;
  wire mux_439_nl;
  wire mux_438_nl;
  wire and_1757_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_2_nl;
  wire[3:0] nor_569_nl;
  wire[3:0] nor_570_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_5_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_2_nl;
  wire and_2681_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_3_nl;
  wire and_2682_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_mux_1_nl;
  wire and_2683_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl;
  wire and_2684_nl;
  wire[7:0] acc_4_nl;
  wire[8:0] nl_acc_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_6_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_or_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_8_nl;
  wire[7:0] acc_5_nl;
  wire[8:0] nl_acc_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_8_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_10_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_11_nl;
  wire[6:0] acc_6_nl;
  wire[7:0] nl_acc_6_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_13_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_14_nl;
  wire[7:0] acc_7_nl;
  wire[8:0] nl_acc_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_22_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_4_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_24_nl;
  wire[7:0] acc_8_nl;
  wire[8:0] nl_acc_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_26_nl;
  wire[7:0] acc_9_nl;
  wire[8:0] nl_acc_9_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl;
  wire[1:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_1_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl;
  wire[7:0] acc_10_nl;
  wire[8:0] nl_acc_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_8_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_28_nl;
  wire[7:0] acc_11_nl;
  wire[8:0] nl_acc_11_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_12_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl;
  wire[4:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl;
  wire[7:0] acc_12_nl;
  wire[8:0] nl_acc_12_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_13_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl;
  wire[4:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl;
  wire i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl;
  wire[3:0] i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl;
  wire[7:0] acc_14_nl;
  wire[8:0] nl_acc_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_5_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_or_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_22_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_8_nl;
  wire[7:0] acc_15_nl;
  wire[8:0] nl_acc_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_4_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_23_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_3_nl;
  wire[7:0] acc_16_nl;
  wire[8:0] nl_acc_16_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_14_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl;
  wire[4:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl;
  wire[7:0] acc_18_nl;
  wire[8:0] nl_acc_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_8_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_15_nl;
  wire and_2685_nl;
  wire[7:0] acc_19_nl;
  wire[8:0] nl_acc_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_25_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_26_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_27_nl;
  wire[7:0] acc_20_nl;
  wire[8:0] nl_acc_20_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl;
  wire[7:0] acc_21_nl;
  wire[8:0] nl_acc_21_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_9_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl;
  wire[4:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl;
  wire[7:0] acc_22_nl;
  wire[8:0] nl_acc_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_29_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_31_nl;
  wire[7:0] acc_23_nl;
  wire[8:0] nl_acc_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_32_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_33_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_34_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_36_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_37_nl;
  wire[7:0] acc_25_nl;
  wire[8:0] nl_acc_25_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl;
  wire[3:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl;
  wire[7:0] acc_26_nl;
  wire[8:0] nl_acc_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_38_nl;
  wire[5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_39_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_40_nl;
  wire[7:0] acc_27_nl;
  wire[8:0] nl_acc_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_25_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_26_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_27_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_28_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_3_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_4_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_5_nl;
  wire[12:0] acc_31_nl;
  wire[13:0] nl_acc_31_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_29_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_30_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_31_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_8_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_32_nl;
  wire[12:0] acc_32_nl;
  wire[13:0] nl_acc_32_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_16_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_18_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_19_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_1_nl;
  wire[12:0] acc_33_nl;
  wire[13:0] nl_acc_33_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_22_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_23_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_9_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_3_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_11_nl;
  wire not_2701_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_24_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_25_nl;
  wire[12:0] acc_34_nl;
  wire[13:0] nl_acc_34_nl;
  wire[10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_13_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_10_nl;
  wire not_2703_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_14_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_15_nl;
  wire[12:0] acc_35_nl;
  wire[13:0] nl_acc_35_nl;
  wire[10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_16_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_12_nl;
  wire not_2705_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_17_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_18_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_7_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_8_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_9_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_10_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_11_nl;
  wire[1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_12_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_13_nl;
  wire[11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_15_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_16_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_17_nl;
  wire[1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_18_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_19_nl;
  wire[11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_20_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_21_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_22_nl;
  wire[1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_23_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_24_nl;
  wire[11:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_25_nl;
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_26_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_27_nl;
  wire[1:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_28_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_29_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_3_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_39_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_1_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_1_nl;

  // Interconnect Declarations for Component Instantiations 
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_28_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_28_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_3_lpi_1_dfm[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]),
      MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_9_nl
      , MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_28_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_42_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_43_nl;
  wire [4:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_42_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_43_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[3:0]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_42_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_43_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_28_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & ac_float_cctor_operator_return_29_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_28_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_64_lpi_1_dfm[3:0]), (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[3:0]),
      ac_float_cctor_operator_return_29_sva);
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_9_nl
      , MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_28_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_4_nl;
  wire [4:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg[3:0]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_10_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_31_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & ac_float_cctor_operator_return_3_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_31_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_65_lpi_1_dfm[3:0]), (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[3:0]),
      ac_float_cctor_operator_return_3_sva);
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_10_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_31_nl};
  wire [12:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0};
  wire [3:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]),
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1, MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0[0])};
  wire [3:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[3:0]),
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1, MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[0])};
  wire [3:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]),
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1, MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl;
  wire [4:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[4]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[3:0]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_7_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_11_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_34_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & ac_float_cctor_operator_return_30_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_34_nl
      = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[3:0]), ac_float_cctor_operator_return_30_sva);
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_11_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_34_nl};
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0};
  wire [3:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]),
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2, MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0[0])};
  wire [3:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]),
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2, MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [3:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]),
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2, MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_10_nl;
  wire [4:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_10_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[3:0]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_10_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_37_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & ac_float_cctor_operator_return_31_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_37_nl
      = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[3:0]),
      ac_float_cctor_operator_return_31_sva);
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_12_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_37_nl};
  wire [12:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0[0])};
  wire [3:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]),
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1[0])};
  wire [3:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]),
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl;
  wire [4:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_12_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[4]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[3:0]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_13_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_13_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_40_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & ac_float_cctor_operator_return_32_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_40_nl
      = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[3:0]),
      ac_float_cctor_operator_return_32_sva);
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_13_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_40_nl};
  wire [12:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0[0])};
  wire [3:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0,
      MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1[0])};
  wire [3:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0,
      MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_16_nl;
  wire [4:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_16_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[3:0]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_16_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_14_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_43_nl;
  wire [5:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_14_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[0])
      & ac_float_cctor_operator_return_42_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_43_nl
      = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2,
      ac_float_cctor_operator_return_42_sva);
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_14_nl
      , MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_43_nl};
  wire [12:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0[0])};
  wire [3:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0,
      MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1[0])};
  wire [3:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0,
      MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_18_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl;
  wire [4:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_18_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_19_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_15_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_46_nl;
  wire [5:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_15_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[0])
      & ac_float_cctor_operator_return_59_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_46_nl
      = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[3:0]),
      ac_float_cctor_operator_return_59_sva);
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_15_nl
      , MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_46_nl};
  wire [12:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[0])};
  wire [3:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0,
      MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva[0])};
  wire [3:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0,
      MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_22_nl;
  wire [4:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_22_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[3:0]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_22_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_28_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_28_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva[3:0]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva);
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_9_nl
      , MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_28_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_45_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_46_nl;
  wire [4:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_45_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_46_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[3:0]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_45_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_46_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_28_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_28_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva);
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      , MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_28_nl};
  wire [12:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva[0])};
  wire [3:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[3:0]),
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1, MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2,
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2,
      (MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl;
  wire [4:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg[3:0]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_3_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_4_nl;
  wire [4:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_3_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[3:0]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl;
  wire [4:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg[4]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg[3:0]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_7_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_7_nl;
  wire [4:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg[4]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_7_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg[3:0]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_7_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_nl;
  wire [4:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg[3:0]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_10_nl;
  wire [4:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_9_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_10_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg[3:0]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_10_nl};
  wire [12:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva[0])};
  wire [3:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[3:0]),
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1, MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire [12:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0};
  wire [3:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]),
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1, MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl;
  wire [4:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg[4]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg[3:0]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_13_nl;
  wire [4:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_12_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg[4]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_13_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg[3:0]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_13_nl};
  wire [12:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva[0])};
  wire [3:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0,
      MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva[0])};
  wire [3:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0,
      MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_13_nl;
  wire [4:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_12_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg[4]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_13_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg[3:0]), MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_13_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl;
  wire [4:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[3:0]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_15_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_16_nl;
  wire [4:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_15_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_16_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[3:0]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_16_nl};
  wire [12:0] nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva[0])};
  wire [3:0] nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0,
      MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva[0])};
  wire [3:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0,
      MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_15_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_16_nl;
  wire [4:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_15_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_16_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[3:0]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_16_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_18_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl;
  wire [4:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_18_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_18_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_19_nl;
  wire [4:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_18_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_19_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_19_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_18_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_19_nl;
  wire [4:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_18_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_19_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_19_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl;
  wire [4:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[3:0]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_21_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_22_nl;
  wire [4:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_21_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_22_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[3:0]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_22_nl};
  wire [12:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva[0])};
  wire [3:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0,
      MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0};
  wire [3:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0,
      MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_21_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_22_nl;
  wire [4:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_21_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_22_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[3:0]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6);
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_mux_22_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_42_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_nl;
  wire [4:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_42_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1,
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[3:0]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_42_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_45_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_nl;
  wire [4:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_45_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[3:0]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_45_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_nl};
  wire [12:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva[0])};
  wire [3:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]),
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1, MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_3_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_4_nl;
  wire [4:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_3_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg[3:0]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_14_lpi_1_dfm[3:0]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva);
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_nl};
  wire [12:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva[0])};
  wire [3:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1,
      MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_6_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_7_nl;
  wire [4:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg[4]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_7_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg[3:0]), MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_7_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_19_lpi_1_dfm[3:0]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva);
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_nl};
  wire [12:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0};
  wire [3:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0,
      MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_9_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_10_nl;
  wire [4:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_9_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_10_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg[3:0]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_mux_10_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_nl
      = MUX_v_4_2_2((operator_ac_float_cctor_e_29_lpi_1_dfm[3:0]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva);
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_nl};
  wire [12:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , 1'b0};
  wire[4:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_57_nl;
  wire [4:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[4:0]),
      ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1}),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_57_nl = ~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = MUX_v_5_2_2(5'b00000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_57_nl);
  wire [11:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      , MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [11:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0};
  wire [11:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0
      , 1'b0};
  wire [11:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1};
  wire [11:0] nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      , MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [11:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0};
  wire [11:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0};
  wire [11:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1
      , 1'b0};
  wire [4:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1};
  wire [11:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0
      , 1'b0};
  wire [4:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      , MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm , operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1};
  wire [4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s;
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s
      = {1'b0, operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_8_nl
      , MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
      , MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s;
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s
      = {1'b0, MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & ac_float_cctor_operator_return_48_sva;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_and_8_nl
      , MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0};
  wire [4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg_s;
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_8_nl
      , MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0};
  wire [4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_10_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_10_nl
      , MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
      , MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0};
  wire [4:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s;
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s
      = {1'b0, MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_10_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva;
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_10_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0};
  wire [4:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_11_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_11_nl
      , MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1};
  wire [4:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s;
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s
      = {1'b0, operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_11_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva;
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_11_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0};
  wire [4:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_12_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_12_nl
      , MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm , operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2};
  wire [4:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s;
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s
      = {1'b0, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_12_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva;
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_12_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0};
  wire [4:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_13_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_and_13_nl
      , MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm , MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [4:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s;
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s
      = {1'b0, MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_13_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva;
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_13_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0};
  wire [4:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_14_nl;
  wire [5:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_14_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva;
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_14_nl
      , MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm , operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1};
  wire [4:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_15_nl;
  wire [5:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_15_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva;
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_and_15_nl
      , MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm , operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1};
  wire [4:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s;
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s
      = {1'b0, operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1};
  wire [12:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0
      , 1'b0};
  wire [4:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      , MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [12:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
      , 1'b0};
  wire [4:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      , MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0};
  wire [12:0] nl_MAC_16_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_16_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0};
  wire [12:0] nl_MAC_15_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_15_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0};
  wire [12:0] nl_MAC_9_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_9_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[0])};
  wire [12:0] nl_MAC_9_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_9_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0};
  wire [12:0] nl_MAC_8_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_8_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0[0])};
  wire [12:0] nl_MAC_8_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_8_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva[0])};
  wire [12:0] nl_MAC_7_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_7_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0[0])};
  wire [12:0] nl_MAC_7_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_7_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva[0])};
  wire [12:0] nl_MAC_6_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_6_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0[0])};
  wire [12:0] nl_MAC_6_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_6_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva[0])};
  wire [12:0] nl_MAC_5_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_5_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0[0])};
  wire [12:0] nl_MAC_5_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_5_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva[0])};
  wire [12:0] nl_MAC_4_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_4_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0[0])};
  wire [12:0] nl_MAC_4_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_4_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva[0])};
  wire [12:0] nl_MAC_3_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_3_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0[0])};
  wire [12:0] nl_MAC_3_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_3_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva[0])};
  wire [12:0] nl_MAC_2_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_2_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[0])};
  wire [12:0] nl_MAC_2_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_2_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_11
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva[0])};
  wire [12:0] nl_MAC_16_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_16_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1[0])};
  wire [12:0] nl_MAC_15_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_15_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1[0])};
  wire [12:0] nl_MAC_14_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_14_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1[0])};
  wire [12:0] nl_MAC_14_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_14_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0};
  wire [12:0] nl_MAC_13_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_13_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_13_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_13_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0};
  wire [12:0] nl_MAC_12_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_12_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[0])};
  wire [12:0] nl_MAC_12_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_12_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva[0])};
  wire [12:0] nl_MAC_11_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_11_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_11_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_11_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva[0])};
  wire [12:0] nl_MAC_10_leading_sign_13_1_1_0_1_rg_mantissa;
  assign nl_MAC_10_leading_sign_13_1_1_0_1_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva[0])};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_3_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_3_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
      , 1'b0};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_2_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_2_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2
      , 1'b0};
  wire [12:0] nl_MAC_2_leading_sign_13_1_1_0_2_rg_mantissa;
  assign nl_MAC_2_leading_sign_13_1_1_0_2_rg_mantissa = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_10_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_29_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_31_nl;
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_nl = MUX_v_5_2_2((signext_5_4(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4:1])),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_10_nl = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_29_nl = MUX_v_2_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1[5:4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_31_nl = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2,
      and_2241_cse);
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_10_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_29_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_31_nl , 1'b0};
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_1_nl;
  wire mux_571_nl;
  wire or_1152_nl;
  wire nor_813_nl;
  wire [4:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_1_nl = MUX_v_5_2_2(z_out_31, ({z_out_32_4
      , z_out_32_3_0}), and_2241_cse);
  assign or_1152_nl = (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | and_2241_cse;
  assign nor_813_nl = ~(MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | and_2241_cse);
  assign mux_571_nl = MUX_s_1_2_2(or_1152_nl, nor_813_nl, MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = MUX_v_5_2_2(5'b00000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_mux_1_nl, mux_571_nl);
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_2_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_19_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_27_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_22_nl;
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_2_nl = MUX_v_5_2_2((signext_5_4(operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0[4:1])),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_19_nl = MUX_s_1_2_2((operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0[0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_27_nl = MUX_v_2_2_2(operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[5:4]),
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_22_nl = MUX_v_4_2_2(operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[3:0]),
      and_2241_cse);
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_2_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_19_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_27_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_22_nl , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_3_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_53_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_54_nl;
  wire mux_572_nl;
  wire or_1153_nl;
  wire nor_815_nl;
  wire [4:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[4]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_3_nl = MUX_s_1_2_2(z_out_32_4, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_53_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5]))
      & and_2241_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_54_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5])
      & and_2241_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_nl
      = MUX1HOT_v_4_3_2(z_out_32_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, {(~ and_2241_cse)
      , operator_13_2_true_AC_TRN_AC_WRAP_1_and_53_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_54_nl});
  assign or_1153_nl = (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | and_2241_cse;
  assign nor_815_nl = ~(MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | and_2241_cse);
  assign mux_572_nl = MUX_s_1_2_2(or_1153_nl, nor_815_nl, MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = MUX_v_5_2_2(5'b00000,
      ({operator_13_2_true_AC_TRN_AC_WRAP_1_mux_3_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_nl}),
      mux_572_nl);
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_4_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_20_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_28_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_23_nl;
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_4_nl = MUX_v_5_2_2((signext_5_4(operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0[4:1])),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_20_nl = MUX_s_1_2_2((operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0[0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_28_nl = MUX_v_2_2_2(operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1,
      and_2241_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_23_nl = MUX_v_4_2_2(operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2,
      and_2241_cse);
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_4_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_20_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_28_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_23_nl , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_5_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_14_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_22_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_20_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_72_nl;
  wire [4:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[4]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl & (~
      MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_5_nl = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_4,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl,
      and_2241_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_20_nl =
      MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_72_nl = ~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_22_nl
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_20_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_72_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_14_nl = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_22_nl,
      and_2241_cse);
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_5_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_14_nl};
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1
      , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_1_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_25_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_20_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_70_nl;
  wire [4:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_4 &
      (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_1_nl = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_itm[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl,
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_70_nl = ~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_20_nl
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_70_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_25_nl = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_itm[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_20_nl,
      and_2317_cse);
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_mux_1_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_25_nl};
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_18_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_23_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_24_nl;
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl = MUX_v_5_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6[5:1]),
      and_2317_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_18_nl = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6[0]),
      and_2317_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_23_nl = MUX_v_2_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4,
      and_2317_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_24_nl = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0,
      and_2317_cse);
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_18_nl , operator_13_2_true_AC_TRN_AC_WRAP_mux_23_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_24_nl , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_3_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_26_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_19_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_69_nl;
  wire [4:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_4 &
      (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_3_nl = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_itm[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl,
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_69_nl = ~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_19_nl
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_69_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_26_nl = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_itm[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_19_nl,
      and_2317_cse);
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_mux_3_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_26_nl};
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
      , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_5_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_27_nl;
  wire[3:0] ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_21_nl;
  wire ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_71_nl;
  wire [4:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_4 &
      (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_5_nl = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_itm[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl,
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_71_nl = ~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_21_nl
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_71_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_27_nl = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_itm[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_21_nl,
      and_2317_cse);
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_mux_5_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_27_nl};
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_6_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_20_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_28_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_29_nl;
  wire [12:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_6_nl = MUX_v_5_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0,
      and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_20_nl = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6,
      and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_28_nl = MUX_v_2_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[5:4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4,
      and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_29_nl = MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0,
      and_2326_cse);
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_mux_6_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_20_nl , operator_13_2_true_AC_TRN_AC_WRAP_mux_28_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_29_nl , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_7_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_14_nl;
  wire [4:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_7_nl = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0, and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_14_nl = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1, and_2326_cse);
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_mux_7_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_14_nl};
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
      , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_9_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_mux_16_nl;
  wire [4:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_9_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0, and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_16_nl = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1, and_2326_cse);
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_mux_9_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_16_nl};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_6_nl;
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_6_nl = MUX_s_1_2_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0]), and_1893_cse);
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_6_nl};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_3_nl;
  wire [3:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_nl
      = ~(MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | and_1893_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_nl = (MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ and_1893_cse)) | (MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_1893_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_3_nl = (~ MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_1893_cse;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]),
      {operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_or_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_3_nl});
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl;
  wire [12:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl
      = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[0]) & (~ and_2438_cse);
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_1_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl;
  wire [3:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_1_nl
      = ~(MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | and_2438_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_nl = (MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ and_2438_cse)) | (MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1
      & and_2438_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl = (~ MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1)
      & and_2438_cse;
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]),
      {operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_1_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_nl});
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_1_nl;
  wire [12:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_1_nl
      = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0[0]) & (~ and_2438_cse);
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2
      , operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_and_1_nl};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_2_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_or_1_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_nl;
  wire [3:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_2_nl
      = ~(MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | and_2438_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_1_nl = (MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ and_2438_cse)) | (MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      & and_2438_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_nl = (~ MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_2438_cse;
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]),
      {operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_nor_2_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_or_1_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_nl});
  wire operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl_1;
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl_1 = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[0]), and_1893_cse);
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_mux_2_nl_1};
  wire operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_nor_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_nl;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_3_nl;
  wire [3:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_nor_nl
      = ~(MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | and_1893_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_nl = (MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ and_1893_cse)) | (MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_1893_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_3_nl = (~ MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_1893_cse;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[3:0]),
      {operator_13_2_true_AC_TRN_AC_WRAP_operator_13_2_true_AC_TRN_AC_WRAP_nor_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_or_nl , operator_13_2_true_AC_TRN_AC_WRAP_and_3_nl});
  wire [12:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])};
  wire [11:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0
      , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_7_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_16_nl;
  wire [4:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_7_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4, and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_16_nl = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0,
      and_2326_cse);
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_7_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_16_nl};
  wire [11:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1
      , 1'b0};
  wire operator_13_2_true_AC_TRN_AC_WRAP_1_mux_9_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_1_mux_18_nl;
  wire [4:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_9_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0,
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4, and_dcpl_2475);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_mux_18_nl = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1,
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, and_dcpl_2475);
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {operator_13_2_true_AC_TRN_AC_WRAP_1_mux_9_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_1_mux_18_nl};
  wire[4:0] operator_13_2_true_AC_TRN_AC_WRAP_2_mux_nl;
  wire[1:0] operator_13_2_true_AC_TRN_AC_WRAP_2_mux_4_nl;
  wire[3:0] operator_13_2_true_AC_TRN_AC_WRAP_2_mux_5_nl;
  wire [11:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a;
  assign operator_13_2_true_AC_TRN_AC_WRAP_2_mux_nl = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6,
      and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_2_mux_4_nl = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4,
      and_2326_cse);
  assign operator_13_2_true_AC_TRN_AC_WRAP_2_mux_5_nl = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0,
      and_2326_cse);
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_2_mux_nl
      , operator_13_2_true_AC_TRN_AC_WRAP_2_mux_4_nl , operator_13_2_true_AC_TRN_AC_WRAP_2_mux_5_nl
      , 1'b0};
  wire [4:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s = {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd11)) input_real_m_rsci (
      .dat(input_real_m_rsc_dat),
      .idat(input_real_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd5)) input_real_e_rsci (
      .dat(input_real_e_rsc_dat),
      .idat(input_real_e_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd11)) input_imag_m_rsci (
      .dat(input_imag_m_rsc_dat),
      .idat(input_imag_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd5)) input_imag_e_rsci (
      .dat(input_imag_e_rsc_dat),
      .idat(input_imag_e_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd5),
  .width(32'sd176)) taps_real_m_rsci (
      .dat(taps_real_m_rsc_dat),
      .idat(taps_real_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd6),
  .width(32'sd80)) taps_real_e_rsci (
      .dat(taps_real_e_rsc_dat),
      .idat(taps_real_e_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd176)) taps_imag_m_rsci (
      .dat(taps_imag_m_rsc_dat),
      .idat(taps_imag_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd80)) taps_imag_e_rsci (
      .dat(taps_imag_e_rsc_dat),
      .idat(taps_imag_e_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd9),
  .width(32'sd11)) return_real_m_rsci (
      .idat(return_real_m_rsci_idat),
      .dat(return_real_m_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd10),
  .width(32'sd5)) return_real_e_rsci (
      .idat(return_real_e_rsci_idat),
      .dat(return_real_e_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd11),
  .width(32'sd11)) return_imag_m_rsci (
      .idat(return_imag_m_rsci_idat),
      .dat(return_imag_m_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd12),
  .width(32'sd5)) return_imag_e_rsci (
      .idat(return_imag_e_rsci_idat),
      .dat(return_imag_e_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_real_m_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(input_real_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_real_e_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(input_real_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_imag_m_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(input_imag_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_imag_e_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(input_imag_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_real_m_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(taps_real_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_real_e_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(taps_real_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_imag_m_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(taps_imag_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_imag_e_triosy_obj (
      .ld(reg_taps_imag_e_triosy_obj_ld_cse),
      .lz(taps_imag_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_real_m_triosy_obj (
      .ld(reg_return_imag_e_triosy_obj_ld_cse),
      .lz(return_real_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_real_e_triosy_obj (
      .ld(reg_return_imag_e_triosy_obj_ld_cse),
      .lz(return_real_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_imag_m_triosy_obj (
      .ld(reg_return_imag_e_triosy_obj_ld_cse),
      .lz(return_imag_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_imag_e_triosy_obj (
      .ld(reg_return_imag_e_triosy_obj_ld_cse),
      .lz(return_imag_e_triosy_lz)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[4:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[4:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_s[3:0]),
      .z(MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[4:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_mx0w2)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_mx0w1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_mx0w1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s[4:0]),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva),
      .s(nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s[4:0]),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva),
      .s(nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_rg_s[4:0]),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva),
      .s(nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva),
      .s(nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s[4:0]),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva),
      .s(nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva),
      .s(nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s[4:0]),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva),
      .s(nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva),
      .s(nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s[4:0]),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva),
      .s(nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva),
      .s(nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_rg_s[4:0]),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva),
      .s(nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva),
      .s(nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[5:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva),
      .s(nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_rg_s[4:0]),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_16_sva_1)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_mx0w0)
    );
  leading_sign_13_1_1_0  MAC_16_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_16_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_70),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_105)
    );
  leading_sign_13_1_1_0  MAC_15_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_15_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_71),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_106)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_72),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_107)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_73),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_108)
    );
  leading_sign_13_1_1_0  MAC_9_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_9_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_74),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_109)
    );
  leading_sign_13_1_1_0  MAC_9_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_9_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_75),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_110)
    );
  leading_sign_13_1_1_0  MAC_8_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_8_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_76),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_111)
    );
  leading_sign_13_1_1_0  MAC_8_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_8_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_77),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_112)
    );
  leading_sign_13_1_1_0  MAC_7_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_7_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_78),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_113)
    );
  leading_sign_13_1_1_0  MAC_7_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_7_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_79),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_114)
    );
  leading_sign_13_1_1_0  MAC_6_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_6_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_80),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_115)
    );
  leading_sign_13_1_1_0  MAC_6_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_6_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_81),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_116)
    );
  leading_sign_13_1_1_0  MAC_5_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_5_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_82),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_117)
    );
  leading_sign_13_1_1_0  MAC_5_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_5_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_83),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_118)
    );
  leading_sign_13_1_1_0  MAC_4_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_4_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_84),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_119)
    );
  leading_sign_13_1_1_0  MAC_4_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_4_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_85),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_120)
    );
  leading_sign_13_1_1_0  MAC_3_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_3_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_86),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_121)
    );
  leading_sign_13_1_1_0  MAC_3_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_3_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_87),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_122)
    );
  leading_sign_13_1_1_0  MAC_2_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_2_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_88),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_123)
    );
  leading_sign_13_1_1_0  MAC_2_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_2_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_89),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_124)
    );
  leading_sign_13_1_1_0  MAC_16_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_16_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_90),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_125)
    );
  leading_sign_13_1_1_0  MAC_15_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_15_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_91),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_126)
    );
  leading_sign_13_1_1_0  MAC_14_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_14_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_92),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_127)
    );
  leading_sign_13_1_1_0  MAC_14_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_14_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_93),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_128)
    );
  leading_sign_13_1_1_0  MAC_13_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_13_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_94),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_129)
    );
  leading_sign_13_1_1_0  MAC_13_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_13_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_95),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_130)
    );
  leading_sign_13_1_1_0  MAC_12_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_12_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_96),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_131)
    );
  leading_sign_13_1_1_0  MAC_12_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_12_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_97),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_132)
    );
  leading_sign_13_1_1_0  MAC_11_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_11_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_98),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_133)
    );
  leading_sign_13_1_1_0  MAC_11_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_11_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_99),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_134)
    );
  leading_sign_13_1_1_0  MAC_10_leading_sign_13_1_1_0_1_rg (
      .mantissa(nl_MAC_10_leading_sign_13_1_1_0_1_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_100),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_135)
    );
  leading_sign_13_1_1_0  MAC_10_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_10_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_101),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_136)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_3_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_3_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_102),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_137)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_2_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_2_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_103),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_138)
    );
  leading_sign_13_1_1_0  MAC_2_leading_sign_13_1_1_0_2_rg (
      .mantissa(nl_MAC_2_leading_sign_13_1_1_0_2_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_104),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_139)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[12:0]),
      .s(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_42)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[12:0]),
      .s(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_43)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[12:0]),
      .s(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_44)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(z_out_45)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(z_out_46)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(z_out_47)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(z_out_48)
    );
  mgc_shift_r_v5 #(.width_a(32'sd13),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[12:0]),
      .s(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_s[4:0]),
      .z(z_out_49)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(z_out_50)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_s[3:0]),
      .z(z_out_51)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_s[3:0]),
      .z(z_out_52)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_a[12:0]),
      .s(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_rg_s[3:0]),
      .z(z_out_53)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_54)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_55)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_56)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_57)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_58)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_59)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_60)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_61)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_62)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_63)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_64)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_rg_a[12:0]),
      .s(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0),
      .z(z_out_65)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_66)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_rg_a[12:0]),
      .s(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0),
      .z(z_out_67)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_68)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_69)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_a[11:0]),
      .s(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_rg_s[4:0]),
      .z(z_out_70)
    );
  fir_core_wait_dp fir_core_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_or_cse =
      and_dcpl_186 | and_dcpl_189;
  assign nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = conv_s2s_5_6(delay_lane_real_e_4_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[29:25]);
  assign MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:0];
  assign nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb
      = ~(MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp | MAC_15_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp);
  assign nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_29_sva);
  assign nl_MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_60_sva);
  assign nl_MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_61_sva);
  assign nl_MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_62_sva);
  assign nl_MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_63_sva);
  assign nl_MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_12_sva);
  assign nl_MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_17_sva);
  assign nl_MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_42_sva);
  assign nl_MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_48_sva);
  assign nl_MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_3_sva);
  assign nl_MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_30_sva);
  assign nl_MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_31_sva);
  assign nl_MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_32_sva);
  assign nl_MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_operator_return_59_sva);
  assign nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb
      = ~(MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign or_1011_tmp = (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & and_dcpl_192) | (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & and_dcpl_199) | (and_dcpl_209 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb))
      | (and_dcpl_1425 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb))
      | (and_dcpl_1427 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb))
      | (and_dcpl_1428 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb))
      | (and_dcpl_1429 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb))
      | (and_dcpl_1430 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb))
      | (and_dcpl_1431 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb))
      | (and_dcpl_1432 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb))
      | (and_dcpl_1433 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb))
      | (and_dcpl_1434 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb))
      | (and_dcpl_1435 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb))
      | (and_dcpl_1436 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb))
      | (and_dcpl_1437 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb))
      | (and_dcpl_1438 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb))
      | (and_dcpl_1439 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb))
      | (and_dcpl_1440 & (~ result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb));
  assign nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = conv_s2s_5_6(delay_lane_imag_e_3_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[24:20]);
  assign MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:0];
  assign nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = conv_s2s_5_6(delay_lane_real_e_3_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[24:20]);
  assign MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = nl_MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:0];
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = conv_s2s_5_6(delay_lane_real_e_8_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:0];
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = conv_s2s_5_6(delay_lane_imag_e_8_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:0];
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = conv_s2s_5_6(delay_lane_real_e_8_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:0];
  assign nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm = conv_s2s_5_6(delay_lane_imag_e_9_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[54:50]);
  assign MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm = nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[5:0];
  assign nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = conv_s2s_5_6(delay_lane_real_e_9_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[54:50]);
  assign MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_5_nl
      = ~((~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_16_nl
      = ~(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm
      = MUX1HOT_v_7_3_2(z_out_7, 7'b1110000, MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_16_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2])});
  assign or_4_nl = (fsm_output[5:3]!=3'b000);
  assign mux_8_cse = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), or_4_nl);
  assign or_6_cse = (fsm_output[5:4]!=2'b00);
  assign MAC_10_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1,
      MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm
      = conv_s2s_6_7(MAC_10_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm =
      nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6:0];
  assign MAC_11_r_ac_float_2_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4,
      MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign MAC_11_r_ac_float_2_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0,
      MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm
      = conv_s2s_6_7({MAC_11_r_ac_float_2_else_and_nl , MAC_11_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm =
      nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6:0];
  assign MAC_12_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0,
      MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm
      = conv_s2s_6_7(MAC_12_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm =
      nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6:0];
  assign MAC_13_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0,
      MAC_13_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm
      = conv_s2s_6_7(MAC_13_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm =
      nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6:0];
  assign MAC_14_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1,
      MAC_14_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm
      = conv_s2s_6_7(MAC_14_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm =
      nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_6_nl
      = ~((~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_17_nl
      = ~(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm
      = MUX1HOT_v_7_3_2(z_out_8, 7'b1110000, MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_17_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2])});
  assign nor_551_m1c = ~(or_dcpl_526 | or_dcpl_527);
  assign or_1078_cse = (fsm_output[3]) | (fsm_output[1]);
  assign and_2663_cse = (fsm_output[3]) & (fsm_output[1]);
  assign mux_536_cse = MUX_s_1_2_2(and_2663_cse, (fsm_output[3]), fsm_output[0]);
  assign or_1077_nl = (fsm_output[3]) | (~ (fsm_output[1]));
  assign mux_535_nl = MUX_s_1_2_2(or_1078_cse, or_1077_nl, fsm_output[0]);
  assign mux_537_nl = MUX_s_1_2_2(mux_536_cse, mux_535_nl, fsm_output[2]);
  assign nor_cse = ~(mux_537_nl | (fsm_output[6:4]!=3'b000));
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_7_nl
      = ~((~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_18_nl
      = ~(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm
      = MUX1HOT_v_7_3_2(z_out_10, 7'b1110000, MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_18_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2])});
  assign nor_552_m1c = ~(or_dcpl_528 | or_dcpl_529);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_1_nl
      = ~((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_19_nl
      = ~(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm
      = MUX1HOT_v_7_3_2((z_out_33[6:0]), 7'b1110000, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_19_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2])});
  assign nor_553_m1c = ~(or_dcpl_530 | or_dcpl_531);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_16_nl
      = ~(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_3
      = MUX_v_7_2_2(z_out_11, 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_16_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_9_nl
      = ~(MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs |
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_37_nl = MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_54_itm = MUX1HOT_v_7_3_2(z_out_9,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_17_nl
      = ~(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_3
      = MUX_v_7_2_2(z_out_12, 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_17_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2}) + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_9_nl
      = ~(ac_float_cctor_operator_return_29_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_37_nl = ac_float_cctor_operator_return_29_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_57_itm = MUX1HOT_v_7_3_2(z_out_4,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_18_nl
      = ~(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_3
      = MUX_v_7_2_2(z_out_18, 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_18_nl);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2}) + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_10_nl
      = ~(ac_float_cctor_operator_return_3_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_41_nl = ac_float_cctor_operator_return_3_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_60_itm = MUX1HOT_v_7_3_2(z_out_19,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign nor_554_m1c = ~(or_dcpl_532 | or_dcpl_533);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_1_nl
      = ~((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_19_nl
      = ~(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_3
      = MUX1HOT_v_7_3_2((z_out_34[6:0]), 7'b1110000, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_19_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2])});
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2}) + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_11_nl
      = ~(ac_float_cctor_operator_return_30_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_45_nl = ac_float_cctor_operator_return_30_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_63_itm = MUX1HOT_v_7_3_2(z_out_22,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign nor_555_m1c = ~(or_dcpl_534 | or_dcpl_535);
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_2_nl
      = ~((~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_20_nl
      = ~(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_3
      = MUX1HOT_v_7_3_2((z_out_35[6:0]), 7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_20_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2])});
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_12_nl
      = ~(ac_float_cctor_operator_return_31_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_49_nl = ac_float_cctor_operator_return_31_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_66_itm = MUX1HOT_v_7_3_2(z_out_5,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign nor_556_m1c = ~(or_dcpl_536 | or_dcpl_537);
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_3_nl
      = ~((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_21_nl
      = ~(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_3
      = MUX1HOT_v_7_3_2((z_out_36[6:0]), 7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_21_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2])});
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_13_nl
      = ~(ac_float_cctor_operator_return_32_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_53_nl = ac_float_cctor_operator_return_32_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_69_itm = MUX1HOT_v_7_3_2(z_out_26,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_4_nl
      = ~((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_22_nl
      = ~(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_3
      = MUX1HOT_v_7_3_2((z_out_37[6:0]), 7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_22_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2])});
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_14_nl
      = ~(ac_float_cctor_operator_return_42_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_57_nl = ac_float_cctor_operator_return_42_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_72_itm = MUX1HOT_v_7_3_2(z_out_23,
      7'b1110000, MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_57_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_16_nl
      = ~(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_3
      = MUX_v_7_2_2(z_out_16, 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_16_nl);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_15_nl
      = ~(ac_float_cctor_operator_return_59_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_61_nl = ac_float_cctor_operator_return_59_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_35_itm = MUX1HOT_v_7_3_2(z_out_15,
      7'b1110000, MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_61_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_17_nl
      = ~(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_3
      = MUX_v_7_2_2(z_out_21, 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_17_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_9_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_37_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_38_itm = MUX1HOT_v_7_3_2(z_out_8,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_7_nl
      = ~((~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_18_nl
      = ~(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_3
      = MUX1HOT_v_7_3_2(z_out_25, 7'b1110000, MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_18_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2])});
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_41_itm = MUX1HOT_v_7_3_2(z_out_27,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg)}) +
      7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_1_nl
      = ~((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_19_nl
      = ~(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_3
      = MUX1HOT_v_7_3_2(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl,
      7'b1110000, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_19_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2])});
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_44_itm = MUX1HOT_v_7_3_2(z_out_14,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg)}) +
      7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_2_nl
      = ~((~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_20_nl
      = ~(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_3
      = MUX1HOT_v_7_3_2(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl,
      7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_20_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2])});
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_47_itm = MUX1HOT_v_7_3_2(z_out_7,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg)}) +
      7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_3_nl
      = ~((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_21_nl
      = ~(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_3
      = MUX1HOT_v_7_3_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl,
      7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_21_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2])});
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_50_itm = MUX1HOT_v_7_3_2(z_out_25,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg)}) +
      7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_4_nl
      = ~((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_22_nl
      = ~(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_3
      = MUX1HOT_v_7_3_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl,
      7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_22_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2])});
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_53_itm = MUX1HOT_v_7_3_2(z_out_10,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg)}) +
      7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_2_nl
      = ~((~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_20_nl
      = ~(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm
      = MUX1HOT_v_7_3_2(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_20_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2])});
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg)}) +
      7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_3_nl
      = ~((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_21_nl
      = ~(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm
      = MUX1HOT_v_7_3_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_21_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2])});
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg)}) +
      7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_4_nl
      = ~((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_22_nl
      = ~(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm
      = MUX1HOT_v_7_3_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_22_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_4_nl
      = ~(and_dcpl_1952 & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2])
      | (fsm_output[4]))) & and_dcpl_2 & and_dcpl_1885)));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_4_nl
      = ~((MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[4]) | and_dcpl_1952);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_23_nl
      = MUX_v_4_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1,
      and_dcpl_1952);
  assign nl_acc_17_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_4_nl})
      + conv_s2u_7_8({(~ and_dcpl_1952) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_23_nl
      , 1'b1});
  assign acc_17_nl = nl_acc_17_nl[7:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl
      = ~(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm
      = MUX_v_7_2_2((readslicef_8_7_1(acc_17_nl)), 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_3_nl
      = ~(and_dcpl_1892 & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2])
      | (fsm_output[4]))) & and_dcpl_2 & and_dcpl_1885)));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_3_nl
      = ~((MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[4]) | and_dcpl_1892);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_21_nl
      = MUX_v_4_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1,
      and_dcpl_1892);
  assign nl_acc_13_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_3_nl})
      + conv_s2u_7_8({(~ and_dcpl_1892) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_21_nl
      , 1'b1});
  assign acc_13_nl = nl_acc_13_nl[7:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl
      = ~(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm
      = MUX_v_7_2_2((readslicef_8_7_1(acc_13_nl)), 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc = and_dcpl_186
      | and_dcpl_243 | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_mx0c2
      | and_dcpl_192;
  assign nor_478_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp[5:4]!=2'b00));
  assign and_1628_cse = (fsm_output[1:0]==2'b11);
  assign or_730_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[5:4]!=2'b01);
  assign nor_479_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5:4]!=2'b00));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse = (~
      and_dcpl_189) & and_dcpl_243;
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_15_nl
      = ~((~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_23_nl
      = ~(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_30_nl
      = MUX1HOT_v_7_3_2(z_out_20, 7'b1110000, MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_23_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_15_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva[21]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_30_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_15_nl);
  assign nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt
      = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1[11:1])
      + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_3_0});
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt
      = nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_ssc = and_dcpl_245
      | and_dcpl_243 | and_dcpl_248 | and_dcpl_251 | and_dcpl_192;
  assign nor_557_m1c = ~(or_dcpl_538 | or_dcpl_539);
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_nl
      = ~((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_24_nl
      = ~(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_nl
      = MUX1HOT_v_7_3_2(z_out_15, 7'b1110000, MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_24_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_nl);
  assign nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt
      = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1[11:1])
      + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0});
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt
      = nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_1_ssc =
      and_dcpl_245 | and_dcpl_243 | and_dcpl_254 | and_dcpl_257 | and_dcpl_192;
  assign nor_558_m1c = ~(or_dcpl_540 | or_dcpl_541);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_14_nl
      = ~((~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_25_nl
      = ~(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_28_nl
      = MUX1HOT_v_7_3_2(z_out_9, 7'b1110000, MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_25_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_14_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva[21]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_28_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_14_nl);
  assign nor_81_cse = ~(ac_float_cctor_operator_return_62_sva | (~ (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign nor_502_nl = ~((MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[6])));
  assign mux_505_nl = MUX_s_1_2_2(nor_502_nl, (fsm_output[6]), MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nor_504_nl = ~((~(ac_float_cctor_operator_return_29_sva | (~ (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_506_nl = MUX_s_1_2_2(mux_505_nl, nor_504_nl, fsm_output[3]);
  assign and_1630_nl = (fsm_output[3]) & (~((~(ac_float_cctor_operator_return_60_sva
      | (~ (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6])));
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, and_1630_nl, fsm_output[2]);
  assign nor_505_nl = ~((~(ac_float_cctor_operator_return_17_sva | (~ (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_506_nl = ~((~(ac_float_cctor_operator_return_48_sva | (~ (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_503_nl = MUX_s_1_2_2(nor_505_nl, nor_506_nl, fsm_output[3]);
  assign nor_507_nl = ~((~(ac_float_cctor_operator_return_42_sva | (~ (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_508_nl = ~((~(ac_float_cctor_operator_return_3_sva | (~ (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_502_nl = MUX_s_1_2_2(nor_507_nl, nor_508_nl, fsm_output[3]);
  assign mux_504_nl = MUX_s_1_2_2(mux_503_nl, mux_502_nl, fsm_output[2]);
  assign mux_508_nl = MUX_s_1_2_2(mux_507_nl, mux_504_nl, fsm_output[5]);
  assign nor_509_nl = ~((~(ac_float_cctor_operator_return_61_sva | (~ (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_510_nl = ~((~(ac_float_cctor_operator_return_63_sva | (~ (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_499_nl = MUX_s_1_2_2(nor_509_nl, nor_510_nl, fsm_output[3]);
  assign nor_511_nl = ~(nor_81_cse | (fsm_output[6]));
  assign nor_512_nl = ~((~(ac_float_cctor_operator_return_12_sva | (~ (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_498_nl = MUX_s_1_2_2(nor_511_nl, nor_512_nl, fsm_output[3]);
  assign mux_500_nl = MUX_s_1_2_2(mux_499_nl, mux_498_nl, fsm_output[2]);
  assign nor_513_nl = ~((~(ac_float_cctor_operator_return_30_sva | (~ (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_514_nl = ~((~(ac_float_cctor_operator_return_32_sva | (~ (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_496_nl = MUX_s_1_2_2(nor_513_nl, nor_514_nl, fsm_output[3]);
  assign nor_515_nl = ~((~(ac_float_cctor_operator_return_31_sva | (~ (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_516_nl = ~((~(ac_float_cctor_operator_return_59_sva | (~ (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_495_nl = MUX_s_1_2_2(nor_515_nl, nor_516_nl, fsm_output[3]);
  assign mux_497_nl = MUX_s_1_2_2(mux_496_nl, mux_495_nl, fsm_output[2]);
  assign mux_501_nl = MUX_s_1_2_2(mux_500_nl, mux_497_nl, fsm_output[5]);
  assign mux_509_nl = MUX_s_1_2_2(mux_508_nl, mux_501_nl, fsm_output[4]);
  assign and_1501_m1c = mux_509_nl & (~(or_tmp_131 | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp));
  assign nor_75_cse = ~(ac_float_cctor_operator_return_61_sva | (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign or_985_cse = and_dcpl_1565 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      | (~ ac_float_cctor_operator_return_60_sva);
  assign or_986_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6;
  assign or_991_cse = and_dcpl_1550 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm);
  assign and_1482_m1c = (((MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_2_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_2_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign and_1486_m1c = and_dcpl_206 & ((~ (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_2_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_2_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign and_1492_m1c = and_dcpl_206 & ((~ (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_59_sva) & nor_137_cse & (~ MAC_11_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp)
      & and_dcpl_164;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_itm = ((~
      or_986_cse) & and_1482_m1c) | ((~ or_985_cse) & and_1486_m1c) | ((~ or_991_cse)
      & and_1492_m1c) | (and_dcpl_1579 & and_1501_m1c);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_3_itm =
      or_986_cse & and_1482_m1c;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_5_itm =
      or_985_cse & and_1486_m1c;
  assign or_761_nl = ac_float_cctor_operator_return_60_sva | (~ nor_tmp_29);
  assign mux_485_nl = MUX_s_1_2_2(mux_tmp_477, or_761_nl, fsm_output[3]);
  assign mux_484_nl = MUX_s_1_2_2((~ mux_tmp_477), (fsm_output[1]), fsm_output[3]);
  assign mux_486_nl = MUX_s_1_2_2((~ mux_485_nl), mux_484_nl, MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp);
  assign and_1488_itm = mux_486_nl & and_dcpl_206 & and_dcpl_633;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_7_itm =
      or_991_cse & and_1492_m1c;
  assign or_765_nl = ac_float_cctor_operator_return_61_sva | (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[4]);
  assign or_764_nl = (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[4]);
  assign mux_490_nl = MUX_s_1_2_2(or_765_nl, or_764_nl, ac_float_cctor_operator_return_30_sva);
  assign mux_491_nl = MUX_s_1_2_2(mux_490_nl, mux_tmp_483, nor_81_cse);
  assign mux_492_nl = MUX_s_1_2_2(mux_491_nl, mux_tmp_483, MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp);
  assign and_1494_itm = (~ mux_492_nl) & and_dcpl_2 & and_dcpl_164;
  assign nor_501_cse = ~((fsm_output[6]) | (fsm_output[3]));
  assign nor_498_nl = ~(ac_float_cctor_operator_return_30_sva | (~ (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[0]) | (~ and_1593_cse));
  assign nor_499_nl = ~((fsm_output[0]) | (~ and_1593_cse));
  assign mux_493_nl = MUX_s_1_2_2(nor_498_nl, nor_499_nl, MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp);
  assign nor_500_nl = ~(ac_float_cctor_operator_return_30_sva | nor_75_cse | (~ (fsm_output[0]))
      | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]));
  assign mux_494_nl = MUX_s_1_2_2(mux_493_nl, nor_500_nl, fsm_output[2]);
  assign and_1496_itm = mux_494_nl & nor_501_cse;
  assign and_1499_itm = (((MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_29_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1090;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_itm = (~
      and_dcpl_1579) & and_1501_m1c;
  assign and_1504_itm = (((MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_61_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1082;
  assign and_1507_itm = (((MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_63_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1090;
  assign and_1510_itm = (((MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_12_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1078;
  assign and_1513_itm = (((MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_17_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1098;
  assign and_1516_itm = (((MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_42_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1102;
  assign and_1519_itm = (((MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_48_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1106;
  assign and_1522_itm = (((MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_3_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1110;
  assign and_1525_itm = (((MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_31_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1102;
  assign and_1528_itm = (((MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_32_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1106;
  assign and_1531_itm = (((MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_59_sva)) | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1110;
  assign and_1534_itm = (((MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_167 & and_dcpl_1082;
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg)}) +
      7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_1_nl
      = ~((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      = ~(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm
      = MUX1HOT_v_7_3_2(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2])});
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg)}) +
      7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      = ~((~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      = ~(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm
      = MUX1HOT_v_7_3_2(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2])});
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg)}) +
      7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      = ~((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      = ~(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm
      = MUX1HOT_v_7_3_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2])});
  assign nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_mx0w0[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1});
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_1_ssc = and_dcpl_186
      | and_dcpl_243 | and_dcpl_209 | and_dcpl_192;
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_nl
      = ~((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_23_nl
      = ~(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_nl
      = MUX1HOT_v_7_3_2(z_out_23, 7'b1110000, MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_23_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_ssc = and_dcpl_186 | and_dcpl_243
      | and_dcpl_209 | and_dcpl_192 | and_dcpl_215;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_1_or_ssc = and_dcpl_186 | and_dcpl_260
      | and_dcpl_209 | and_dcpl_198;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_5_nl
      = ~(and_dcpl_2029 & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2])
      | (fsm_output[4]))) & and_dcpl_2 & and_dcpl_1885)));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_5_nl
      = ~((MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[4]) | and_dcpl_2029);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_24_nl
      = MUX_v_4_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1,
      and_dcpl_2029);
  assign nl_acc_24_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_5_nl})
      + conv_s2u_7_8({(~ and_dcpl_2029) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_24_nl
      , 1'b1});
  assign acc_24_nl = nl_acc_24_nl[7:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl
      = ~(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm
      = MUX_v_7_2_2((readslicef_8_7_1(acc_24_nl)), 7'b1110000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl);
  assign nor_559_m1c = ~(or_dcpl_543 | or_dcpl_544);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg)}) +
      7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      = ~((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      = ~(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm
      = MUX1HOT_v_7_3_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2])});
  assign nor_560_m1c = ~(or_dcpl_546 | or_dcpl_548);
  assign nor_561_m1c = ~(or_dcpl_550 | or_dcpl_552);
  assign MAC_13_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0,
      MAC_13_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm
      = conv_s2s_6_7(MAC_13_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm =
      nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6:0];
  assign nor_562_m1c = ~(or_dcpl_554 | or_dcpl_555);
  assign MAC_14_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1,
      MAC_14_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm
      = conv_s2s_6_7(MAC_14_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm =
      nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6:0];
  assign and_269_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2])
      & nor_98_cse;
  assign and_272_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2])))
      & nor_98_cse;
  assign and_275_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[1]);
  assign and_278_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1[1])));
  assign mux_197_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_1078_cse);
  assign mux_195_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, and_1628_cse);
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, mux_tmp_188, fsm_output[3]);
  assign mux_198_nl = MUX_s_1_2_2(mux_197_nl, mux_196_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_2_ssc = and_dcpl_186
      | (~(mux_198_nl | (fsm_output[6]))) | and_dcpl_192;
  assign and_568_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2])
      & nor_98_cse;
  assign and_571_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2])))
      & nor_98_cse;
  assign and_574_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign and_577_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1[1])));
  assign nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2});
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign or_361_cse = (fsm_output[3]) | (fsm_output[0]);
  assign mux_204_nl = MUX_s_1_2_2(not_tmp_212, nor_tmp_6, or_1078_cse);
  assign mux_575_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, and_1628_cse);
  assign mux_203_nl = MUX_s_1_2_2(mux_575_nl, nor_tmp_6, fsm_output[3]);
  assign mux_205_nl = MUX_s_1_2_2(mux_204_nl, mux_203_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_3_ssc = and_dcpl_186
      | (~(mux_205_nl | (fsm_output[6]))) | and_dcpl_192;
  assign and_618_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2])
      & nor_98_cse;
  assign and_621_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2])))
      & nor_98_cse;
  assign and_624_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign and_627_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1[1])));
  assign nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1});
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign mux_213_nl = MUX_s_1_2_2(not_tmp_307, nor_tmp_6, fsm_output[3]);
  assign mux_211_nl = MUX_s_1_2_2(mux_tmp_147, mux_tmp_65, fsm_output[0]);
  assign mux_212_nl = MUX_s_1_2_2(mux_211_nl, nor_tmp_6, fsm_output[3]);
  assign mux_214_nl = MUX_s_1_2_2(mux_213_nl, mux_212_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_4_ssc = and_dcpl_186
      | (~(mux_214_nl | (fsm_output[6]))) | and_dcpl_192;
  assign and_705_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2])
      & nor_98_cse;
  assign and_708_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2])))
      & nor_98_cse;
  assign and_711_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[1]);
  assign and_714_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1[1])));
  assign nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2});
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign mux_220_nl = MUX_s_1_2_2(not_tmp_307, and_1593_cse, fsm_output[3]);
  assign mux_219_nl = MUX_s_1_2_2(not_tmp_284, nor_tmp_6, fsm_output[3]);
  assign mux_221_nl = MUX_s_1_2_2(mux_220_nl, mux_219_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_5_ssc = and_dcpl_186
      | (~(mux_221_nl | (fsm_output[6]))) | and_dcpl_192;
  assign and_784_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2])
      & nor_98_cse;
  assign and_787_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2])))
      & nor_98_cse;
  assign and_790_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[1]);
  assign and_793_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1[1])));
  assign nor_235_nl = ~((fsm_output[3]) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]));
  assign mux_225_nl = MUX_s_1_2_2(not_tmp_284, and_1593_cse, fsm_output[3]);
  assign mux_226_nl = MUX_s_1_2_2(nor_235_nl, mux_225_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_6_ssc = and_dcpl_186
      | (~(mux_226_nl | (fsm_output[6]))) | and_dcpl_192;
  assign and_870_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2])
      & nor_98_cse;
  assign and_873_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2])))
      & nor_98_cse;
  assign and_876_itm = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[1]);
  assign and_879_itm = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1[1])));
  assign nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2});
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_7_ssc = and_dcpl_186
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1
      | and_dcpl_192;
  assign and_1318_itm = nor_469_cse & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2])
      & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1;
  assign and_1321_itm = nor_469_cse & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2])))
      & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1;
  assign and_1324_itm = and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1])
      & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1;
  assign and_1327_itm = and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1])))
      & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1;
  assign MAC_9_r_ac_float_1_else_and_nl = operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1
      & MAC_9_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  assign MAC_9_r_ac_float_1_else_and_1_nl = MUX_v_5_2_2(5'b00000, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2,
      MAC_9_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm =
      conv_s2s_6_7({MAC_9_r_ac_float_1_else_and_nl , MAC_9_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_ssc = ~(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva[21]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign or_378_nl = (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]);
  assign mux_234_nl = MUX_s_1_2_2(mux_tmp_223, or_378_nl, fsm_output[2]);
  assign and_362_ssc = (~ mux_234_nl) & and_dcpl_206;
  assign or_972_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_16_tmp[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_8_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_16_tmp[6]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_5_ssc = and_dcpl_243 | and_dcpl_222
      | and_dcpl_192;
  assign nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(z_out_68[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1});
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = conv_s2u_11_12(z_out_69[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1});
  assign MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm =
      nl_MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = (z_out_49[12:1]) + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1});
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = conv_s2u_11_12(z_out_70[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0});
  assign MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm =
      nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_16_sva_1[12:1])
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1});
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = (z_out_48[12:1]) + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0});
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(z_out_69[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1});
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_mx0w1[11:1])
      + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_3_0});
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl =
      ~ MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      = MUX_v_5_2_2(5'b00000, operator_i_m_1_lpi_1_dfm_mx0w3_10_6, result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl =
      ~ MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl
      = MUX_v_6_2_2(6'b000000, operator_i_m_1_lpi_1_dfm_mx0w3_5_0, result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      = MUX_v_5_2_2(5'b00000, operator_i_m_1_lpi_1_dfm_mx0w3_10_6, MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl
      = MUX_v_6_2_2(6'b000000, operator_i_m_1_lpi_1_dfm_mx0w3_5_0, MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = conv_s2u_11_12({result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      , result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl})
      + conv_s2u_11_12({result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      , result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl});
  assign MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm =
      nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_mx0w1[11:1])
      + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_3_0});
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl =
      ~ MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      = MUX_v_5_2_2(5'b00000, operator_r_m_1_lpi_1_dfm_mx0w4_10_6, result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_32_nl);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl =
      ~ MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl
      = MUX_v_6_2_2(6'b000000, operator_r_m_1_lpi_1_dfm_mx0w4_5_0, result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_33_nl);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      = MUX_v_5_2_2(5'b00000, operator_r_m_1_lpi_1_dfm_mx0w4_10_6, MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl
      = MUX_v_6_2_2(6'b000000, operator_r_m_1_lpi_1_dfm_mx0w4_5_0, MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm
      = conv_s2u_11_12({result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      , result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_nl})
      + conv_s2u_11_12({result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      , result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_nl});
  assign MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm =
      nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_8_ssc =
      and_dcpl_243 | and_dcpl_367 | and_dcpl_370 | and_dcpl_192;
  assign MAC_13_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1,
      MAC_13_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm
      = conv_s2s_6_7(MAC_13_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm =
      nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_9_ssc =
      and_dcpl_243 | and_dcpl_373 | and_dcpl_376 | and_dcpl_192;
  assign MAC_14_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1,
      MAC_14_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm
      = conv_s2s_6_7(MAC_14_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm =
      nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_10_ssc
      = and_dcpl_243 | and_dcpl_399 | and_dcpl_402 | and_dcpl_192;
  assign MAC_15_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1,
      MAC_15_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm
      = conv_s2s_6_7(MAC_15_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm =
      nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6:0];
  assign nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (z_out_48[12:1]) + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0});
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_8_ssc = and_dcpl_243
      | and_dcpl_399 | and_dcpl_402 | and_dcpl_194;
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl
      = ~((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      = ~(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_nl
      = MUX1HOT_v_7_3_2(z_out_14, 7'b1110000, MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl);
  assign nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3[11:1])
      + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0});
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(z_out_70[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0});
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = conv_s2u_11_12(z_out_68[11:1]) + conv_s2u_11_12({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0});
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm
      = nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
      | and_dcpl_452 | and_dcpl_455;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1
      | and_dcpl_478 | and_dcpl_481 | and_dcpl_484 | and_dcpl_487 | and_dcpl_198;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_1_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1
      | and_dcpl_521 | and_dcpl_524 | and_dcpl_484 | and_dcpl_487 | and_dcpl_198;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_4_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_212;
  assign and_631_itm = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2])
      & nor_98_cse;
  assign and_634_itm = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2])))
      & nor_98_cse;
  assign and_1610_nl = (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[1]) & (fsm_output[4]);
  assign nor_265_nl = ~((~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | (fsm_output[1]) | (fsm_output[4]));
  assign mux_270_nl = MUX_s_1_2_2(and_1610_nl, nor_265_nl, fsm_output[2]);
  assign and_636_itm = mux_270_nl & and_dcpl_2 & nor_469_cse;
  assign nor_266_nl = ~((MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      | (fsm_output[1]));
  assign mux_271_nl = MUX_s_1_2_2(nor_266_nl, nor_tmp_29, fsm_output[3]);
  assign and_640_itm = mux_271_nl & (~ (fsm_output[6])) & not_tmp_212 & and_dcpl_633;
  assign nor_267_nl = ~((~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[4]));
  assign nor_268_nl = ~((~ (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[0]) | (~ nor_tmp_26));
  assign mux_272_nl = MUX_s_1_2_2(nor_267_nl, nor_268_nl, fsm_output[3]);
  assign and_642_itm = mux_272_nl & and_dcpl_637;
  assign nand_44_nl = ~((fsm_output[3]) & (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ (fsm_output[0])) & and_1593_cse);
  assign or_904_nl = (fsm_output[3]) | (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]);
  assign mux_273_nl = MUX_s_1_2_2(nand_44_nl, or_904_nl, fsm_output[2]);
  assign nor_270_itm = ~(mux_273_nl | (fsm_output[6]));
  assign and_647_itm = and_dcpl_188 & (~ (fsm_output[0])) & (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign or_905_nl = (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[2]) | (~ (fsm_output[6]));
  assign or_906_nl = (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_907_nl = (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_284_nl = MUX_s_1_2_2(or_906_nl, or_907_nl, fsm_output[2]);
  assign mux_285_nl = MUX_s_1_2_2(or_905_nl, mux_284_nl, fsm_output[3]);
  assign or_908_nl = (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_909_nl = (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_282_nl = MUX_s_1_2_2(or_908_nl, or_909_nl, fsm_output[2]);
  assign or_910_nl = (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_911_nl = (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_281_nl = MUX_s_1_2_2(or_910_nl, or_911_nl, fsm_output[2]);
  assign mux_283_nl = MUX_s_1_2_2(mux_282_nl, mux_281_nl, fsm_output[3]);
  assign mux_286_nl = MUX_s_1_2_2(mux_285_nl, mux_283_nl, fsm_output[5]);
  assign or_912_nl = (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_913_nl = (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_278_nl = MUX_s_1_2_2(or_912_nl, or_913_nl, fsm_output[2]);
  assign or_914_nl = (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_915_nl = (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_277_nl = MUX_s_1_2_2(or_914_nl, or_915_nl, fsm_output[2]);
  assign mux_279_nl = MUX_s_1_2_2(mux_278_nl, mux_277_nl, fsm_output[3]);
  assign or_916_nl = (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_917_nl = (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_275_nl = MUX_s_1_2_2(or_916_nl, or_917_nl, fsm_output[2]);
  assign or_918_nl = (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_919_nl = (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_274_nl = MUX_s_1_2_2(or_918_nl, or_919_nl, fsm_output[2]);
  assign mux_276_nl = MUX_s_1_2_2(mux_275_nl, mux_274_nl, fsm_output[3]);
  assign mux_280_nl = MUX_s_1_2_2(mux_279_nl, mux_276_nl, fsm_output[5]);
  assign mux_287_nl = MUX_s_1_2_2(mux_286_nl, mux_280_nl, fsm_output[4]);
  assign nor_286_itm = ~(mux_287_nl | or_tmp_131);
  assign and_652_itm = and_dcpl_647 & (~ (fsm_output[0])) & (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_655_itm = and_dcpl_647 & (~ (fsm_output[0])) & (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign and_660_itm = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign and_663_itm = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_666_itm = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign and_670_itm = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_663;
  assign and_674_itm = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign and_677_itm = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_680_itm = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_663;
  assign and_684_itm = and_dcpl_679 & (~ (fsm_output[0])) & (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_3_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1
      | and_dcpl_689 | and_dcpl_692;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_4_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1
      | and_dcpl_689 | and_dcpl_692;
  assign or_467_cse = (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_5_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1
      | and_dcpl_854 | and_dcpl_857;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_6_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1
      | and_dcpl_854 | and_dcpl_857;
  assign or_987_cse = nor_539_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0;
  assign or_988_cse = nor_540_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_8_ssc = ((~
      or_988_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c1)
      | ((~ or_987_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c2)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_1_ssc = or_988_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_3_ssc = or_987_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_ssc = and_dcpl_189
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c1
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c2
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c3
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c4;
  assign or_981_cse = (~ ac_float_cctor_operator_return_62_sva) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
      | nor_195_cse;
  assign or_982_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6;
  assign and_1587_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]==2'b01);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse =
      MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[4:0]),
      5'b01111, and_1587_cse);
  assign or_983_cse = and_dcpl_1562 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0
      | (~ ac_float_cctor_operator_return_61_sva);
  assign or_984_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6;
  assign or_989_cse = and_dcpl_1568 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_10_ssc = ((~
      or_984_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c1)
      | ((~ or_983_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c2)
      | ((~ or_989_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c4)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c8
      | (and_1587_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c9);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_9_ssc = or_984_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_11_ssc =
      or_983_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_13_ssc =
      or_989_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_14_ssc =
      (~ and_1587_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c9;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_2_ssc = and_dcpl_189
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c1
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c2
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c3
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c4
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c5
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c6
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c7
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c8
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c9
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c10
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c11
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c12
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c13
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c14
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c15
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c16
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c17
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c18
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c19
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c20
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c21
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c22
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c23;
  assign or_993_cse = and_dcpl_1554 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm);
  assign or_994_cse = and_dcpl_1551 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm);
  assign or_979_cse = and_dcpl_1355 | (~ ac_float_cctor_operator_return_63_sva) |
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0;
  assign or_980_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6;
  assign nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb
      = ~(MAC_1_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp | MAC_1_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp);
  assign nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_1_ssc = and_dcpl_189
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_192 | and_dcpl_194 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c5
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c6;
  assign or_977_cse = and_dcpl_1363 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0;
  assign or_978_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6;
  assign or_992_cse = and_dcpl_1565 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign or_975_cse = and_dcpl_1551 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0;
  assign or_976_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6;
  assign or_990_cse = and_dcpl_1562 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_13_ssc = ((~
      or_976_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c1)
      | ((~ or_975_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c2)
      | ((~ or_990_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c4)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c8;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_31_ssc =
      or_976_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_33_ssc =
      or_975_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_35_ssc =
      or_990_cse & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_5_ssc = and_dcpl_189
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c1
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c2
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c3
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c4
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c5
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c6
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c7
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c8;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_8_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1
      | and_dcpl_452 | and_dcpl_455;
  assign or_973_cse = and_dcpl_1547 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0;
  assign or_974_cse = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_cse =
      and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_dcpl_198;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_cse
      = and_dcpl_189 | and_dcpl_209 | and_dcpl_212;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_1_cse
      = and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_dcpl_212;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_2_cse
      = and_dcpl_189 | and_dcpl_209 | and_dcpl_198;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_1_cse = and_dcpl_189
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_194 | and_dcpl_195 | and_dcpl_212;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_3_cse = and_dcpl_189
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_194 | and_dcpl_195 | and_dcpl_198;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_4_cse = and_dcpl_189
      | and_dcpl_209 | and_dcpl_194 | and_dcpl_198;
  assign nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb
      = ~(MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp | MAC_16_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp);
  assign nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm);
  assign nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb
      = ~(MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm);
  assign or_1065_tmp = (and_dcpl_209 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb))
      | (and_dcpl_192 & MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | (and_dcpl_1425 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb))
      | (and_dcpl_1427 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb))
      | (and_dcpl_1428 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb))
      | (and_dcpl_1429 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb))
      | (and_dcpl_1430 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb))
      | (and_dcpl_1431 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb))
      | (and_dcpl_1432 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb))
      | (and_dcpl_1433 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb))
      | (and_dcpl_1434 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb))
      | (and_dcpl_1435 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb))
      | (and_dcpl_1436 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb))
      | (and_dcpl_1437 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb))
      | (and_dcpl_1438 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb))
      | (and_dcpl_1439 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb))
      | (and_dcpl_1440 & (~ result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb));
  assign or_967_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5:4]!=2'b01);
  assign or_900_cse = (fsm_output[1]) | (fsm_output[4]);
  assign or_968_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5:4]!=2'b01);
  assign or_966_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5:4]!=2'b01);
  assign and_969_rgt = and_dcpl_964 & and_dcpl_963;
  assign or_486_nl = (or_966_cse & (fsm_output[0])) | (fsm_output[1]);
  assign mux_353_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_486_nl);
  assign mux_354_nl = MUX_s_1_2_2(not_tmp_307, mux_353_nl, fsm_output[3]);
  assign mux_355_nl = MUX_s_1_2_2(mux_354_nl, mux_tmp_149, fsm_output[2]);
  assign or_487_rgt = mux_355_nl | (fsm_output[6]);
  assign nor_137_cse = ~((fsm_output[1:0]!=2'b00));
  assign and_1593_cse = (fsm_output[1]) & (fsm_output[4]) & (fsm_output[5]);
  assign nor_138_nl = ~(nor_137_cse | (fsm_output[5:4]!=2'b00));
  assign mux_80_cse = MUX_s_1_2_2(nor_138_nl, nor_tmp_6, fsm_output[3]);
  assign and_1331_rgt = and_dcpl_1142 & and_dcpl_1267;
  assign mux_395_nl = MUX_s_1_2_2(not_tmp_307, mux_tmp_65, fsm_output[3]);
  assign mux_396_nl = MUX_s_1_2_2(mux_395_nl, mux_80_cse, fsm_output[2]);
  assign nor_53_nl = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0!=2'b01));
  assign mux_400_nl = MUX_s_1_2_2(mux_tmp_393, mux_396_nl, nor_53_nl);
  assign or_590_rgt = mux_400_nl | (fsm_output[6]);
  assign nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_21_ssc = or_590_rgt & (~ and_dcpl_192);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_11_ssc = ((~(mux_tmp_393 | (fsm_output[6])))
      | and_dcpl_192) & (and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_1331_rgt
      | or_590_rgt);
  assign nor_469_cse = ~((fsm_output[3]) | (fsm_output[0]));
  assign and_462_ssc = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2])
      & nor_98_cse;
  assign and_465_ssc = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2])))
      & nor_98_cse;
  assign and_468_ssc = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign and_471_ssc = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1])));
  assign mux_448_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), or_1078_cse);
  assign or_707_nl = (~ (fsm_output[0])) | (~ (fsm_output[1])) | (fsm_output[4]);
  assign mux_447_nl = MUX_s_1_2_2(or_707_nl, (fsm_output[4]), fsm_output[3]);
  assign mux_449_nl = MUX_s_1_2_2(mux_448_nl, mux_447_nl, fsm_output[2]);
  assign mux_245_nl = MUX_s_1_2_2(or_tmp_154, or_tmp_153, fsm_output[3]);
  assign or_392_nl = (fsm_output[4:3]!=2'b01);
  assign mux_246_nl = MUX_s_1_2_2(mux_245_nl, or_392_nl, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_7_ssc = (((~ mux_449_nl) & and_dcpl_2)
      | and_dcpl_192) & (~((~ mux_246_nl) & and_dcpl_2));
  assign and_506_ssc = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2])
      & nor_98_cse;
  assign and_509_ssc = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2])))
      & nor_98_cse;
  assign and_512_ssc = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign and_515_ssc = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1])));
  assign mux_453_nl = MUX_s_1_2_2((~ or_900_cse), (fsm_output[4]), fsm_output[3]);
  assign mux_451_nl = MUX_s_1_2_2(or_tmp_154, mux_tmp_247, fsm_output[0]);
  assign mux_452_nl = MUX_s_1_2_2(mux_451_nl, (fsm_output[4]), fsm_output[3]);
  assign mux_454_nl = MUX_s_1_2_2(mux_453_nl, mux_452_nl, fsm_output[2]);
  assign mux_250_nl = MUX_s_1_2_2((~ (fsm_output[4])), or_tmp_153, fsm_output[3]);
  assign mux_249_nl = MUX_s_1_2_2(or_tmp_154, (fsm_output[4]), fsm_output[3]);
  assign mux_251_nl = MUX_s_1_2_2(mux_250_nl, mux_249_nl, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_8_ssc = (((~ mux_454_nl) & and_dcpl_2)
      | and_dcpl_192) & (~((~ mux_251_nl) & and_dcpl_2));
  assign and_581_ssc = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2])
      & nor_98_cse;
  assign and_584_ssc = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2])))
      & nor_98_cse;
  assign and_587_ssc = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign and_590_ssc = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1])));
  assign nor_205_nl = ~((fsm_output[3]) | (fsm_output[1]) | (fsm_output[4]));
  assign mux_463_nl = MUX_s_1_2_2(nor_205_nl, mux_tmp_257, fsm_output[2]);
  assign or_399_nl = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[4]);
  assign mux_264_nl = MUX_s_1_2_2((fsm_output[4]), or_399_nl, fsm_output[3]);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, (~ mux_tmp_257), fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_10_ssc = (((~ mux_463_nl) & and_dcpl_2)
      | and_dcpl_192) & (~(mux_265_nl & and_dcpl_2));
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_8_cse = and_dcpl_209 | and_dcpl_198;
  assign nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = (z_out_49[12:1]) + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1});
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt
      = nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_6_ssc
      = and_dcpl_361 | and_dcpl_364 | and_dcpl_1575 | and_dcpl_1578 | and_dcpl_420
      | and_dcpl_423 | and_dcpl_194;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_7_ssc
      = and_dcpl_432 | and_dcpl_435 | and_dcpl_1575 | and_dcpl_1578 | and_dcpl_194;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_8_cse
      = and_dcpl_199 | and_dcpl_194;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0 = $signed((input_real_m_rsci_idat))
      * $signed((taps_real_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0 = $signed((input_imag_m_rsci_idat))
      * $signed((taps_imag_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0 = $signed((input_real_m_rsci_idat))
      * $signed((taps_imag_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0 = $signed((input_imag_m_rsci_idat))
      * $signed((taps_real_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0 = $signed(delay_lane_real_m_0_sva)
      * $signed((taps_real_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0 = $signed(delay_lane_imag_m_0_sva)
      * $signed((taps_imag_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0 = $signed(delay_lane_real_m_0_sva)
      * $signed((taps_imag_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0 = $signed(delay_lane_imag_m_0_sva)
      * $signed((taps_real_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0 = $signed(delay_lane_real_m_1_sva)
      * $signed((taps_real_m_rsci_idat[32:22]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0 = $signed(delay_lane_imag_m_1_sva)
      * $signed((taps_imag_m_rsci_idat[32:22]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0 = $signed(delay_lane_real_m_1_sva)
      * $signed((taps_imag_m_rsci_idat[32:22]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0 = $signed(delay_lane_imag_m_1_sva)
      * $signed((taps_real_m_rsci_idat[32:22]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0 = $signed(delay_lane_real_m_2_sva)
      * $signed((taps_real_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0 = $signed(delay_lane_imag_m_2_sva)
      * $signed((taps_imag_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0 = $signed(delay_lane_real_m_2_sva)
      * $signed((taps_imag_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0 = $signed(delay_lane_imag_m_2_sva)
      * $signed((taps_real_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0 = $signed(delay_lane_real_m_3_sva)
      * $signed((taps_real_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0 = $signed(delay_lane_imag_m_3_sva)
      * $signed((taps_imag_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0 = $signed(delay_lane_real_m_3_sva)
      * $signed((taps_imag_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0 = $signed(delay_lane_imag_m_3_sva)
      * $signed((taps_real_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0 = $signed(delay_lane_real_m_4_sva)
      * $signed((taps_real_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0 = $signed(delay_lane_imag_m_4_sva)
      * $signed((taps_imag_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0 = $signed(delay_lane_real_m_4_sva)
      * $signed((taps_imag_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0 = $signed(delay_lane_imag_m_4_sva)
      * $signed((taps_real_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0 = $signed(delay_lane_real_m_5_sva)
      * $signed((taps_real_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0 = $signed(delay_lane_imag_m_5_sva)
      * $signed((taps_imag_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0 = $signed(delay_lane_real_m_5_sva)
      * $signed((taps_imag_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0 = $signed(delay_lane_imag_m_5_sva)
      * $signed((taps_real_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0 = $signed(delay_lane_real_m_6_sva)
      * $signed((taps_real_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0 = $signed(delay_lane_imag_m_6_sva)
      * $signed((taps_imag_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0 = $signed(delay_lane_real_m_6_sva)
      * $signed((taps_imag_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0 = $signed(delay_lane_imag_m_6_sva)
      * $signed((taps_real_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0 = $signed(delay_lane_real_m_13_sva)
      * $signed((taps_real_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0 = $signed(delay_lane_imag_m_13_sva)
      * $signed((taps_imag_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0 = $signed(delay_lane_real_m_14_sva)
      * $signed((taps_real_m_rsci_idat[175:165]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0 = $signed(delay_lane_imag_m_14_sva)
      * $signed((taps_imag_m_rsci_idat[175:165]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0 = $signed(delay_lane_real_m_7_sva)
      * $signed((taps_real_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0 = $signed(delay_lane_imag_m_7_sva)
      * $signed((taps_imag_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0 = $signed(delay_lane_real_m_7_sva)
      * $signed((taps_imag_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0 = $signed(delay_lane_imag_m_7_sva)
      * $signed((taps_real_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0 = $signed(delay_lane_real_m_8_sva)
      * $signed((taps_real_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0 = $signed(delay_lane_imag_m_8_sva)
      * $signed((taps_imag_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0 = $signed(delay_lane_real_m_8_sva)
      * $signed((taps_imag_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0 = $signed(delay_lane_imag_m_8_sva)
      * $signed((taps_real_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0 = $signed(delay_lane_real_m_9_sva)
      * $signed((taps_real_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0 = $signed(delay_lane_imag_m_9_sva)
      * $signed((taps_imag_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0 = $signed(delay_lane_real_m_9_sva)
      * $signed((taps_imag_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0 = $signed(delay_lane_imag_m_9_sva)
      * $signed((taps_real_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0 = $signed(delay_lane_real_m_10_sva)
      * $signed((taps_real_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0 = $signed(delay_lane_imag_m_10_sva)
      * $signed((taps_imag_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0 = $signed(delay_lane_real_m_10_sva)
      * $signed((taps_imag_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0 = $signed(delay_lane_imag_m_10_sva)
      * $signed((taps_real_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0 = $signed(delay_lane_real_m_11_sva)
      * $signed((taps_real_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0 = $signed(delay_lane_imag_m_11_sva)
      * $signed((taps_imag_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0 = $signed(delay_lane_real_m_11_sva)
      * $signed((taps_imag_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0 = $signed(delay_lane_imag_m_11_sva)
      * $signed((taps_real_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0 = $signed(delay_lane_real_m_12_sva)
      * $signed((taps_real_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0 = $signed(delay_lane_imag_m_12_sva)
      * $signed((taps_imag_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0 = $signed(delay_lane_real_m_12_sva)
      * $signed((taps_imag_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0 = $signed(delay_lane_imag_m_12_sva)
      * $signed((taps_real_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0 = $signed(delay_lane_real_m_13_sva)
      * $signed((taps_imag_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0 = $signed(delay_lane_imag_m_13_sva)
      * $signed((taps_real_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0 = $signed(delay_lane_real_m_14_sva)
      * $signed((taps_imag_m_rsci_idat[175:165]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0 = $signed(delay_lane_imag_m_14_sva)
      * $signed((taps_real_m_rsci_idat[175:165]));
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva)
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[5:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva)
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1 = conv_s2s_5_6({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0})
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[5:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1 = conv_s2s_5_6({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1}) +
      6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1[5:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva)
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[5:0];
  assign MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_13_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_28_lpi_1_dfm_mx0);
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva)
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2[5:0];
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_12_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_27_lpi_1_dfm_mx0);
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_10_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_25_lpi_1_dfm_mx0);
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_9_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_24_lpi_1_dfm_mx0);
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_8_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_23_lpi_1_dfm_mx0);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6 = MUX_v_6_2_2(6'b000000,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_11_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_26_lpi_1_dfm_mx0);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_4_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
      or_973_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_5_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
      or_974_cse);
  assign MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_4_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_5_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6 = MUX_v_6_2_2(6'b000000,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_7_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_22_lpi_1_dfm_mx0);
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1 = conv_s2s_5_6(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1 = conv_s2s_5_6(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[5:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[5:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[5:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[5:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1 = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1)
      + 6'b000001;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1 = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[5:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = conv_s2s_5_6({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0})
      + 6'b000001;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:0];
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_28_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0[4:0]),
      or_985_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_29_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0[4:0]),
      or_986_cse);
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_28_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_29_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_40_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
      or_993_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_41_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
      or_994_cse);
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_40_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_41_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_24_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0[4:0]),
      or_983_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_25_nl = MUX_v_5_2_2(5'b01111,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0,
      or_984_cse);
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_24_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_25_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_38_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0[4:0]),
      or_991_cse);
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_38_nl)
      - $signed(operator_ac_float_cctor_e_61_lpi_1_dfm);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_20_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_4_lpi_1_dfm_1_5_0[4:0]),
      or_981_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_21_nl = MUX_v_5_2_2(5'b01111,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_4_lpi_1_dfm_1_4_0,
      or_982_cse);
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_20_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_21_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_36_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0[4:0]),
      or_989_cse);
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_36_nl)
      - $signed(operator_ac_float_cctor_e_62_lpi_1_dfm);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_16_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_5_lpi_1_dfm_1_5_0[4:0]),
      or_979_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_17_nl = MUX_v_5_2_2(5'b01111,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_5_lpi_1_dfm_1_4_0,
      or_980_cse);
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_16_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_17_nl);
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_15_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_30_lpi_1_dfm_mx0);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_12_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_6_lpi_1_dfm_1_5_0[4:0]),
      or_977_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_13_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_6_lpi_1_dfm_1_5_0[4:0]),
      or_978_cse);
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_12_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_13_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_39_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1_5_0[4:0]),
      or_992_cse);
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_39_nl)
      - $signed(operator_ac_float_cctor_e_31_lpi_1_dfm);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_8_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0[4:0]),
      or_975_cse);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_9_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0[4:0]),
      or_976_cse);
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_8_nl)
      - $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_9_nl);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_37_nl = MUX_v_5_2_2(5'b01111,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0[4:0]),
      or_990_cse);
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_37_nl)
      - $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2);
  assign MAC_2_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1,
      MAC_2_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1
      = conv_s2s_6_7(MAC_2_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1[6:0];
  assign MAC_3_r_ac_float_4_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
      & MAC_3_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  assign MAC_3_r_ac_float_4_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1,
      MAC_3_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1
      = conv_s2s_6_7({MAC_3_r_ac_float_4_else_and_nl , MAC_3_r_ac_float_4_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1[6:0];
  assign MAC_4_r_ac_float_4_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0
      & MAC_4_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  assign MAC_4_r_ac_float_4_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1,
      MAC_4_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1
      = conv_s2s_6_7({MAC_4_r_ac_float_4_else_and_nl , MAC_4_r_ac_float_4_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1[6:0];
  assign MAC_5_r_ac_float_4_else_and_nl = MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_5
      & MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  assign MAC_5_r_ac_float_4_else_and_1_nl = MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_4
      & MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  assign MAC_5_r_ac_float_4_else_and_2_nl = MUX_v_4_2_2(4'b0000, MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0,
      MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1
      = conv_s2s_6_7({MAC_5_r_ac_float_4_else_and_nl , MAC_5_r_ac_float_4_else_and_1_nl
      , MAC_5_r_ac_float_4_else_and_2_nl}) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1[6:0];
  assign MAC_3_r_ac_float_2_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0
      & MAC_3_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  assign MAC_3_r_ac_float_2_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1,
      MAC_3_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1
      = conv_s2s_6_7({MAC_3_r_ac_float_2_else_and_nl , MAC_3_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1[6:0];
  assign MAC_4_r_ac_float_2_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0
      & MAC_4_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  assign MAC_4_r_ac_float_2_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1,
      MAC_4_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1
      = conv_s2s_6_7({MAC_4_r_ac_float_2_else_and_nl , MAC_4_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1[6:0];
  assign MAC_5_r_ac_float_2_else_and_nl = operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1
      & MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  assign MAC_5_r_ac_float_2_else_and_1_nl = operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0
      & MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  assign MAC_5_r_ac_float_2_else_and_2_nl = MUX_v_4_2_2(4'b0000, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1,
      MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1
      = conv_s2s_6_7({MAC_5_r_ac_float_2_else_and_nl , MAC_5_r_ac_float_2_else_and_1_nl
      , MAC_5_r_ac_float_2_else_and_2_nl}) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1[6:0];
  assign MAC_6_r_ac_float_2_else_and_nl = MUX_v_2_2_2(2'b00, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1,
      MAC_6_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign MAC_6_r_ac_float_2_else_and_1_nl = MUX_v_4_2_2(4'b0000, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2,
      MAC_6_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1
      = conv_s2s_6_7({MAC_6_r_ac_float_2_else_and_nl , MAC_6_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1[6:0];
  assign MAC_7_r_ac_float_2_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
      MAC_7_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign MAC_7_r_ac_float_2_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
      MAC_7_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1
      = conv_s2s_6_7({MAC_7_r_ac_float_2_else_and_nl , MAC_7_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1[6:0];
  assign MAC_8_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1}),
      MAC_8_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1
      = conv_s2s_6_7(MAC_8_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1[6:0];
  assign MAC_16_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1,
      MAC_16_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1
      = conv_s2s_6_7(MAC_16_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1[6:0];
  assign MAC_2_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1,
      MAC_2_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1
      = conv_s2s_6_7(MAC_2_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1[6:0];
  assign MAC_3_r_ac_float_3_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0
      & MAC_3_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_3_r_ac_float_3_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1,
      MAC_3_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1
      = conv_s2s_6_7({MAC_3_r_ac_float_3_else_and_nl , MAC_3_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1[6:0];
  assign MAC_4_r_ac_float_3_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0
      & MAC_4_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_4_r_ac_float_3_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1,
      MAC_4_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1
      = conv_s2s_6_7({MAC_4_r_ac_float_3_else_and_nl , MAC_4_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1[6:0];
  assign MAC_5_r_ac_float_3_else_and_nl = MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5
      & MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_5_r_ac_float_3_else_and_1_nl = MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      & MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_5_r_ac_float_3_else_and_2_nl = MUX_v_4_2_2(4'b0000, MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0,
      MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1
      = conv_s2s_6_7({MAC_5_r_ac_float_3_else_and_nl , MAC_5_r_ac_float_3_else_and_1_nl
      , MAC_5_r_ac_float_3_else_and_2_nl}) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1[6:0];
  assign MAC_6_r_ac_float_3_else_and_nl = MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5
      & MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_6_r_ac_float_3_else_and_1_nl = MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4
      & MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_6_r_ac_float_3_else_and_2_nl = MUX_v_4_2_2(4'b0000, MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0,
      MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1
      = conv_s2s_6_7({MAC_6_r_ac_float_3_else_and_nl , MAC_6_r_ac_float_3_else_and_1_nl
      , MAC_6_r_ac_float_3_else_and_2_nl}) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1[6:0];
  assign MAC_7_r_ac_float_3_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
      MAC_7_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign MAC_7_r_ac_float_3_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
      MAC_7_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1
      = conv_s2s_6_7({MAC_7_r_ac_float_3_else_and_nl , MAC_7_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1[6:0];
  assign MAC_8_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1}),
      MAC_8_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1
      = conv_s2s_6_7(MAC_8_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1[6:0];
  assign MAC_6_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1,
      MAC_6_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1
      = conv_s2s_6_7(MAC_6_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1[6:0];
  assign MAC_7_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1}),
      MAC_7_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1
      = conv_s2s_6_7(MAC_7_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1[6:0];
  assign MAC_8_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1}),
      MAC_8_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1
      = conv_s2s_6_7(MAC_8_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1[6:0];
  assign MAC_3_r_ac_float_1_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
      & MAC_3_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  assign MAC_3_r_ac_float_1_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1,
      MAC_3_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1
      = conv_s2s_6_7({MAC_3_r_ac_float_1_else_and_nl , MAC_3_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[6:0];
  assign MAC_4_r_ac_float_1_else_and_nl = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
      & MAC_4_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  assign MAC_4_r_ac_float_1_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2,
      MAC_4_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1
      = conv_s2s_6_7({MAC_4_r_ac_float_1_else_and_nl , MAC_4_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[6:0];
  assign MAC_6_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1,
      MAC_6_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1
      = conv_s2s_6_7(MAC_6_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[6:0];
  assign MAC_7_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1}),
      MAC_7_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1
      = conv_s2s_6_7(MAC_7_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[6:0];
  assign MAC_8_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1}),
      MAC_8_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1
      = conv_s2s_6_7(MAC_8_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_54_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_14_lpi_1_dfm_mx0[10]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_55_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_14_lpi_1_dfm_mx0[10])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_14_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_54_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_55_nl});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_18);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_18);
  assign MAC_5_r_ac_float_1_else_and_nl = MUX_v_2_2_2(2'b00, operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0,
      MAC_5_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign MAC_5_r_ac_float_1_else_and_1_nl = MUX_v_4_2_2(4'b0000, operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1,
      MAC_5_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1
      = conv_s2s_6_7({MAC_5_r_ac_float_1_else_and_nl , MAC_5_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[6:0];
  assign MAC_16_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1,
      MAC_16_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1
      = conv_s2s_6_7(MAC_16_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_54_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_55_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_28_ssc
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_22);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_44_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_22);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_19);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_19);
  assign MAC_1_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1,
      MAC_1_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1
      = conv_s2s_6_7(MAC_1_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:0];
  assign MAC_1_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1,
      MAC_1_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1
      = conv_s2s_6_7(MAC_1_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1[6:0];
  assign MAC_1_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1,
      MAC_1_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1
      = conv_s2s_6_7(MAC_1_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1[6:0];
  assign MAC_1_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1,
      MAC_1_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1
      = conv_s2s_6_7(MAC_1_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1[6:0];
  assign MAC_2_r_ac_float_1_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0
      & MAC_2_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm;
  assign MAC_2_r_ac_float_1_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1,
      MAC_2_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1
      = conv_s2s_6_7({MAC_2_r_ac_float_1_else_and_nl , MAC_2_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1[6:0];
  assign MAC_2_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1,
      MAC_2_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1
      = conv_s2s_6_7(MAC_2_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1[6:0];
  assign MAC_15_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1,
      MAC_15_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1
      = conv_s2s_6_7(MAC_15_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1[6:0];
  assign MAC_15_r_ac_float_2_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1,
      MAC_15_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1
      = conv_s2s_6_7(MAC_15_r_ac_float_2_else_and_nl) + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1[6:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1
      =  -(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1
      =  -(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_7_ssc
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4]) | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_15_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24);
  assign operator_r_m_8_lpi_1_dfm_mx0w6_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6, {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_7_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_15_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_86_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_15_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_66_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_86_nl);
  assign operator_r_m_8_lpi_1_dfm_mx0w6_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_66_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_7_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_85_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_15_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_85_nl);
  assign operator_r_m_8_lpi_1_dfm_mx0w6_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_64_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_7_ssc);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1[3:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg) + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1
      =  -(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_2_sva_1[3:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg) + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_2_sva_1[3:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg) + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_8_ssc
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4]) | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_17_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20);
  assign operator_r_m_9_lpi_1_dfm_mx0w6_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6, {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_8_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_17_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_94_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_17_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_94_nl);
  assign operator_r_m_9_lpi_1_dfm_mx0w6_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_8_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_82_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_17_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_68_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_82_nl);
  assign operator_r_m_9_lpi_1_dfm_mx0w6_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_68_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_8_ssc);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_2_sva_1[3:0];
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg) + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_3_sva_1[3:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg) + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_3_sva_1[3:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg) + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_5_ssc
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_32);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_11_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_32);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_3_sva_1[3:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg) + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_16);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_16);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_3_sva_1[3:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg) + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_48_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_48_nl);
  assign operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_17_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_17_nl);
  assign operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_ssc);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_4_sva_1[3:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg) + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_42);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_42);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_4_sva_1[3:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg) + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_6_ssc
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4]) | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_28);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_13_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_28);
  assign operator_r_m_7_lpi_1_dfm_mx0w4_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6, {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_6_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_13_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_28});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_92_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_13_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_92_nl);
  assign operator_r_m_7_lpi_1_dfm_mx0w4_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_6_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_83_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_13_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_65_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_83_nl);
  assign operator_r_m_7_lpi_1_dfm_mx0w4_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_65_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_6_ssc);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_4_sva_1[3:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg) + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_4_sva_1[3:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg) + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6[4]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6[4])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_45_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_45_nl);
  assign operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_34_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_34_nl);
  assign operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_ssc);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_5_sva_1[3:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg) + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_40);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_40);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_5_sva_1[3:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg) + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_5_sva_1[3:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg) + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_5_sva_1[3:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg) + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_42_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_11_lpi_1_dfm_mx0[10]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_43_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_11_lpi_1_dfm_mx0[10])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_11_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_42_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_43_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_62_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_63_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_17);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_17);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_6_sva_1[3:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg) + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1[3:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg) + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1[3:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg) + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_6_sva_1[3:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg) + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_62_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_lpi_1_dfm_mx0[10]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_63_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_lpi_1_dfm_mx0[10])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_62_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_63_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_7_sva_1[3:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg) + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1[3:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg) + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1[3:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg) + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_7_sva_1[3:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg) + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_46_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_12_lpi_1_dfm_mx0[10]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_47_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_12_lpi_1_dfm_mx0[10])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_12_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_46_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_47_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_50_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_51_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_26);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_26);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_8_sva_1[3:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg) + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1[3:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg) + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_8_sva_1[3:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg) + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_8_sva_1[3:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg) + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1[4])})
      + 3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0}) +
      3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0 , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[4])})
      + 3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4})
      + 3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4})
      + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[4])}) + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[5:4])})
      + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4})
      + 3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[4])}) +
      3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0})
      + 3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0})
      + 3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1
      , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[4])}) +
      3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1})
      + 3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0})
      + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1})
      + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0})
      + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[5:4])})
      + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1[5:4])})
      + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1[3:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_15_sva_1[3:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1})
      + 3'b001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1})
      + 3'b001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_50_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_13_lpi_1_dfm_mx0[10]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_51_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_13_lpi_1_dfm_mx0[10])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_13_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_50_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_51_nl});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_26_ssc
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4])
      | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_42_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1[3:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_sva_1[3:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
      , (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[5:4])})
      + 3'b001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0 , (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[5:4])})
      + 3'b001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:0];
  assign my_complex_float_t_cctor_imag_operator_return_4_sva_mx0w1 = ~((operator_r_m_lpi_1_dfm_mx0w6_10_6!=5'b00000)
      | (operator_r_m_lpi_1_dfm_mx0w6_5_4!=2'b00) | (operator_r_m_lpi_1_dfm_mx0w6_3_0!=4'b0000));
  assign my_complex_float_t_cctor_real_operator_return_9_sva_mx0w1 = ~((operator_i_m_9_lpi_1_dfm_mx0w10_10_6!=5'b00000)
      | (operator_i_m_9_lpi_1_dfm_mx0w10_5_4!=2'b00) | (operator_i_m_9_lpi_1_dfm_mx0w10_3_0!=4'b0000));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_operator_return_2_sva_mx0w2 = ~((operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      = ~((operator_i_m_1_lpi_1_dfm_mx0w3_10_6!=5'b00000) | (operator_i_m_1_lpi_1_dfm_mx0w3_5_0!=6'b000000));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp
      = ~((operator_r_m_1_lpi_1_dfm_mx0w4_10_6!=5'b00000) | (operator_r_m_1_lpi_1_dfm_mx0w4_5_0!=6'b000000));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_operator_return_46_sva_mx0w2 = ~((operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign my_complex_float_t_cctor_imag_operator_return_3_sva_mx0w3 = ~((operator_r_m_15_lpi_1_dfm_mx0w4_10_6!=5'b00000)
      | (operator_r_m_15_lpi_1_dfm_mx0w4_5_4!=2'b00) | (operator_r_m_15_lpi_1_dfm_mx0w4_3_0!=4'b0000));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign my_complex_float_t_cctor_imag_operator_return_13_sva_mx0w2 = ~((operator_i_m_6_lpi_1_dfm_mx0w4_10_6!=5'b00000)
      | (operator_i_m_6_lpi_1_dfm_mx0w4_5_4!=2'b00) | (operator_i_m_6_lpi_1_dfm_mx0w4_3_0!=4'b0000));
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign my_complex_float_t_cctor_imag_operator_return_14_sva_mx0w2 = ~((operator_i_m_7_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_i_m_7_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_i_m_7_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_itm_mx0w7
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_100 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[0])));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign my_complex_float_t_cctor_imag_operator_return_sva_mx0w6 = ~((operator_i_m_8_lpi_1_dfm_mx0w10_10_6!=5'b00000)
      | (operator_i_m_8_lpi_1_dfm_mx0w10_5_4!=2'b00) | (operator_i_m_8_lpi_1_dfm_mx0w10_3_0!=4'b0000));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign my_complex_float_t_cctor_real_operator_return_10_sva_mx0w6 = ~((operator_r_m_2_lpi_1_dfm_mx0w6_10_6!=5'b00000)
      | (operator_r_m_2_lpi_1_dfm_mx0w6_5_4!=2'b00) | (operator_r_m_2_lpi_1_dfm_mx0w6_3_0!=4'b0000));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[1:0]))
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign my_complex_float_t_cctor_real_operator_return_11_sva_mx0w5 = ~((operator_r_m_3_lpi_1_dfm_mx0w6_10_6!=5'b00000)
      | (operator_r_m_3_lpi_1_dfm_mx0w6_5_4!=2'b00) | (operator_r_m_3_lpi_1_dfm_mx0w6_3_0!=4'b0000));
  assign my_complex_float_t_cctor_real_operator_return_12_sva_mx0w5 = ~((operator_r_m_4_lpi_1_dfm_mx0w5_10_6!=5'b00000)
      | (operator_r_m_4_lpi_1_dfm_mx0w5_5_4!=2'b00) | (operator_r_m_4_lpi_1_dfm_mx0w5_3_0!=4'b0000));
  assign my_complex_float_t_cctor_real_operator_return_4_sva_mx0w5 = ~((operator_r_m_14_lpi_1_dfm_mx0w5_10_6!=5'b00000)
      | (operator_r_m_14_lpi_1_dfm_mx0w5_5_4!=2'b00) | (operator_r_m_14_lpi_1_dfm_mx0w5_3_0!=4'b0000));
  assign ac_float_cctor_operator_return_12_sva_mx0w1 = ~((operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_operator_return_16_sva_mx0w2 = ~((operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign ac_float_cctor_operator_return_27_sva_mx0w1 = ~((operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_operator_return_17_sva_mx0w2 = ~((operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2)})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_operator_return_42_sva_mx0w1 = ~((operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_operator_return_47_sva_mx0w2 = ~((operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_5_4!=2'b00) | (operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_3_0!=4'b0000));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_operator_return_57_sva_mx0w1 = ~((operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_operator_return_48_sva_mx0w2 = ~((operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_5_4!=2'b00) | (operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_3_0!=4'b0000));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_20_nl
      = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4[0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[4]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_4
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_20_nl &
      (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_27_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_78_nl = ~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_3_0
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_27_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_78_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_58_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_59_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_42_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_11_lpi_1_dfm_mx0[10]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_43_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_11_lpi_1_dfm_mx0[10])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_11_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_42_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_43_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_46_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_12_lpi_1_dfm_mx0[10]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_47_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_12_lpi_1_dfm_mx0[10])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_12_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_46_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_47_nl});
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(({operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_4 , operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_3_0}))
      - $signed(operator_ac_float_cctor_e_21_lpi_1_dfm_mx0);
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_32_nl = MUX_v_5_2_2(5'b01111,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2,
      or_987_cse);
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nand_nl
      = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1[0])
      & or_988_cse);
  assign not_nl = ~ or_988_cse;
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nor_nl
      = ~(MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2,
      4'b1111, not_nl));
  assign nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_mux_32_nl)
      + conv_s2s_5_6({MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nand_nl
      , MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_e_ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_nor_nl})
      + 6'b000001;
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva_1[3:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_10_sva_1[3:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1
      =  -(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_10_sva_1[3:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1
      =  -(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_10_sva_1[3:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_11_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_11_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:11]),
      (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1
      =  -(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_11_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_11_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_12_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_12_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:11]),
      (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1
      =  -(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_12_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_12_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_13_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_13_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:11]),
      (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_13_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_13_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_14_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_14_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:11]),
      (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_14_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_14_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6({operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_4 , operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_3_0})
      + conv_s2s_5_6({(~ operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_4) , (~ operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_3_0)})
      + 6'b000001;
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1
      =  -ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_15_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_15_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1[1]);
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_1_lpi_1_dfm_mx0);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1
      =  -(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:11]),
      (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_58_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_15_lpi_1_dfm_mx0[10]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_59_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_15_lpi_1_dfm_mx0[10])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_15_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_58_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_59_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_54_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_14_lpi_1_dfm_mx0[10]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_55_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_14_lpi_1_dfm_mx0[10])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_14_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_54_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_55_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_50_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_13_lpi_1_dfm_mx0[10]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_51_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_13_lpi_1_dfm_mx0[10])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_13_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_50_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_51_nl});
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva)})
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1})
      + conv_u2s_4_7(operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_15_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_61_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp
      = MUX1HOT_v_7_3_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_61_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nor_521_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4])
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[0]));
  assign or_803_nl = nor_521_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1]);
  assign operator_ac_float_cctor_e_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0,
      or_803_nl);
  assign nor_522_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[4])
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1);
  assign or_804_nl = nor_522_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0;
  assign operator_ac_float_cctor_e_1_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2,
      or_804_nl);
  assign MAC_16_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_1_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_1_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_1_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6[4]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6[4])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_49_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_49_nl);
  assign operator_ac_float_cctor_m_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_18_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_18_nl);
  assign operator_ac_float_cctor_m_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1 = conv_s2s_11_12({(~
      operator_ac_float_cctor_m_1_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_1_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_1_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_62_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_63_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
      | nor_522_cse);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1])
      | nor_521_cse);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva)})
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2})
      + conv_u2s_4_7(operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_14_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_57_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp
      = MUX1HOT_v_7_3_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_57_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_15_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_15_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_15_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nor_523_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0!=2'b00));
  assign or_805_ssc = nor_523_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6;
  assign operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_4 = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0[0])
      & or_805_ssc;
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl = ~ or_805_ssc;
  assign operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_3_0 = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1,
      4'b1111, ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl);
  assign nor_524_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0!=2'b00));
  assign or_806_ssc = nor_524_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0;
  assign operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_4 = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0[0])
      & or_806_ssc;
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_1_nl = ~ or_806_ssc;
  assign operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_3_0 = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      4'b1111, ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_1_nl);
  assign MAC_15_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_35_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_35_lpi_1_dfm_1_5_0!=6'b000000));
  assign MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_20_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_20_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6[4]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6[4])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_35_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_35_nl);
  assign operator_ac_float_cctor_m_20_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_30_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_30_nl);
  assign operator_ac_float_cctor_m_20_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1
      = conv_s2s_11_12({(~ operator_ac_float_cctor_m_35_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_35_lpi_1_dfm_1_5_0)})
      + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_58_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_59_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
      | nor_524_cse);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      | nor_523_cse);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0)})
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_13_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_53_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp
      = MUX1HOT_v_7_3_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_14_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_14_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_14_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_62_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1})
      + conv_u2s_4_7(MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_13_nl
      = ~(MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs |
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_53_nl = MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp
      = MUX1HOT_v_7_3_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_14_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp,
      MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_14_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_14_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva)})
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_12_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_49_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp
      = MUX1HOT_v_7_3_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_13_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_13_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_13_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_61_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1})
      + conv_u2s_4_7(operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_12_nl
      = ~(MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_49_nl = MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp
      = MUX1HOT_v_7_3_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_13_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp,
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_13_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_13_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva)})
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_11_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_45_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp
      = MUX1HOT_v_7_3_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_12_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_12_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_12_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_34_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1})
      + conv_u2s_4_7(operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_11_nl
      = ~(MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs |
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_45_nl = MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp
      = MUX1HOT_v_7_3_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_12_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp,
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_12_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_12_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0)})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_10_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_41_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp
      = MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_11_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_11_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_11_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_33_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_10_nl
      = ~(MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_41_nl = MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp
      = MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_11_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp,
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_11_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_11_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0}) + conv_s2s_6_7({1'b1
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0)})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0}) + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_8_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_33_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_16_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_8_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0)})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_8_nl
      = ~(ac_float_cctor_operator_return_48_sva | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_33_nl = ac_float_cctor_operator_return_48_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_63_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_8_nl
      = ~(MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_33_nl = MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp,
      ac_float_cctor_operator_return_17_sva);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ operator_ac_float_cctor_e_31_lpi_1_dfm)}) + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1})
      + conv_u2s_4_7(operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign MAC_8_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_58_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_58_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_58_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_8_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_43_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_43_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_43_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_30_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6[4]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_31_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6[4])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_58_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_30_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_31_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_39_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_76_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_39_nl);
  assign operator_ac_float_cctor_m_58_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_76_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_26_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_95_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_26_nl);
  assign operator_ac_float_cctor_m_58_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_95_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_8_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_8_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_8_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_812_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6;
  assign operator_ac_float_cctor_e_13_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
      or_812_nl);
  assign or_814_nl = and_dcpl_1550 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      | (~ ac_float_cctor_operator_return_12_sva);
  assign operator_ac_float_cctor_e_28_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
      or_814_nl);
  assign MAC_8_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_28_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_28_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_28_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_13_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_13_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6[4]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6[4])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_50_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_50_nl);
  assign operator_ac_float_cctor_m_13_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_19_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_19_nl);
  assign operator_ac_float_cctor_m_13_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_28_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_28_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_28_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_30_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0[4]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_31_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0[4])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      & ac_float_cctor_operator_return_12_sva) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_8_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_7_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_57_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_57_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_57_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_7_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_42_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_42_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_42_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_26_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6[4]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_27_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6[4])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_57_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_26_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_27_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_40_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_77_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_40_nl);
  assign operator_ac_float_cctor_m_57_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_77_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_27_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_96_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_27_nl);
  assign operator_ac_float_cctor_m_57_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_96_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_820_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6;
  assign operator_ac_float_cctor_e_12_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1_4_0,
      or_820_nl);
  assign or_822_nl = and_dcpl_1554 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      | (~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_ac_float_cctor_e_27_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_7_lpi_1_dfm_1_5_0[4:0]),
      or_822_nl);
  assign MAC_7_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_27_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_27_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_27_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_12_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_12_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6[4]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6[4])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_40_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_40_nl);
  assign operator_ac_float_cctor_m_12_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_20_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_20_nl);
  assign operator_ac_float_cctor_m_12_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_27_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_27_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_27_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_26_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_27_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0[4])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      & MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_7_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1_4_0[4]))));
  assign MAC_6_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_56_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_56_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_56_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_6_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_41_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_41_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_41_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_22_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0[4]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_23_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0[4])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_22_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6[4]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_23_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6[4])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_56_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_22_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_23_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_41_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_93_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_41_nl);
  assign operator_ac_float_cctor_m_56_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_93_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_32_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_97_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_32_nl);
  assign operator_ac_float_cctor_m_56_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_97_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_6_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_6_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_6_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_828_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6;
  assign operator_ac_float_cctor_e_11_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1_4_0,
      or_828_nl);
  assign or_830_nl = and_dcpl_1557 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
      | (~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign operator_ac_float_cctor_e_26_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_6_lpi_1_dfm_1_5_0[4:0]),
      or_830_nl);
  assign MAC_6_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_26_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_26_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_26_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_11_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_11_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6[4]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6[4])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_41_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_41_nl);
  assign operator_ac_float_cctor_m_11_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_21_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_21_nl);
  assign operator_ac_float_cctor_m_11_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_26_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_26_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_26_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_22_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_23_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0[4])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
      & MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_6_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1_4_0[4]))));
  assign MAC_5_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_55_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_55_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_55_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_5_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_40_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_40_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_40_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_18_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0[4]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_19_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0[4])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_18_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6[4]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_19_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6[4])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_55_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_18_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_19_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_42_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_94_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_42_nl);
  assign operator_ac_float_cctor_m_55_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_94_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_33_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_98_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_33_nl);
  assign operator_ac_float_cctor_m_55_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_98_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_18_ssc);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_5_lpi_1_dfm_1_4_0[4]))));
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
      & ac_float_cctor_operator_return_63_sva) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_5_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_836_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6;
  assign operator_ac_float_cctor_e_10_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1_5_0[4:0]),
      or_836_nl);
  assign or_838_nl = and_dcpl_1463 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
      | (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign operator_ac_float_cctor_e_25_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_5_lpi_1_dfm_1_5_0[4:0]),
      or_838_nl);
  assign MAC_5_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_25_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_25_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_25_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_10_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_10_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6[4]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6[4])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_46_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_46_nl);
  assign operator_ac_float_cctor_m_10_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_29_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_29_nl);
  assign operator_ac_float_cctor_m_10_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_25_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_25_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_25_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_18_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_19_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0[4])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
      & MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_5_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_4_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_54_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_54_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_54_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_4_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_39_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_39_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_39_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_14_ssc = (~
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6[4])) & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_15_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6[4])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_39_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_15_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_51_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_100_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_51_nl);
  assign operator_ac_float_cctor_m_39_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_100_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_42_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_103_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_42_nl);
  assign operator_ac_float_cctor_m_39_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_103_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_14_ssc);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_4_lpi_1_dfm_1_4_0[4]))));
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
      & ac_float_cctor_operator_return_62_sva) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_4_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign nor_534_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0);
  assign or_844_nl = nor_534_cse | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6;
  assign operator_ac_float_cctor_e_9_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1_4_0,
      or_844_nl);
  assign or_846_nl = nor_479_cse | (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0;
  assign operator_ac_float_cctor_e_24_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_4_lpi_1_dfm_1_5_0[4:0]),
      or_846_nl);
  assign MAC_4_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_24_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_24_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_24_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_9_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_9_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[4]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[4])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_51_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_51_nl);
  assign operator_ac_float_cctor_m_9_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_22_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_22_nl);
  assign operator_ac_float_cctor_m_9_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_24_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_24_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_24_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
      & MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_4_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1_4_0[4]))));
  assign MAC_3_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_53_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_53_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_53_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_3_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_38_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_38_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_38_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_10_ssc = (~
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4])) & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_11_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6[4])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_38_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_10_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_11_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_56_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_74_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_56_nl);
  assign operator_ac_float_cctor_m_38_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_74_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_26_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_108_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_26_nl);
  assign operator_ac_float_cctor_m_38_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_108_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_10_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6[4]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_11_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6[4])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_53_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_10_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_11_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_36_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_70_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_36_nl);
  assign operator_ac_float_cctor_m_53_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_70_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_20_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_90_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_20_nl);
  assign operator_ac_float_cctor_m_53_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_90_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_10_ssc);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0[4]))));
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0
      & ac_float_cctor_operator_return_61_sva) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign nor_536_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0);
  assign or_852_nl = nor_536_cse | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6;
  assign operator_ac_float_cctor_e_8_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1_4_0,
      or_852_nl);
  assign or_854_nl = nor_199_cse | (~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0;
  assign operator_ac_float_cctor_e_23_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_3_lpi_1_dfm_1_5_0[4:0]),
      or_854_nl);
  assign MAC_3_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_23_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_23_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_23_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_8_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_8_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6[4]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6[4])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_42_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_42_nl);
  assign operator_ac_float_cctor_m_8_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_23_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_23_nl);
  assign operator_ac_float_cctor_m_8_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_23_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_23_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_23_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_10_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_11_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
      & MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) |
      (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_3_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1_4_0[4]))));
  assign MAC_2_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_52_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_52_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_52_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_2_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_37_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_37_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_37_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_6_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_7_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_37_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_6_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_7_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_43_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_102_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_43_nl);
  assign operator_ac_float_cctor_m_37_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_102_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_30_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_99_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_30_nl);
  assign operator_ac_float_cctor_m_37_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_99_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_6_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6[4]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_7_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6[4])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_52_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_6_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_7_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_37_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_73_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_37_nl);
  assign operator_ac_float_cctor_m_52_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_73_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_23_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_91_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_23_nl);
  assign operator_ac_float_cctor_m_52_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_91_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      & ac_float_cctor_operator_return_60_sva) | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_860_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6;
  assign operator_ac_float_cctor_e_7_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_4_0,
      or_860_nl);
  assign or_862_nl = and_dcpl_1568 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
      | (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign operator_ac_float_cctor_e_22_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_2_lpi_1_dfm_1_5_0[4:0]),
      or_862_nl);
  assign MAC_2_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_22_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_22_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_22_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_7_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_7_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_6_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6[4]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_7_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6[4])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_6_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_7_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_43_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_43_nl);
  assign operator_ac_float_cctor_m_7_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_24_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_24_nl);
  assign operator_ac_float_cctor_m_7_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_6_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_22_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_22_lpi_1_dfm_1_5_4)
      , (~ operator_ac_float_cctor_m_22_lpi_1_dfm_1_3_0)}) + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_6_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_7_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
      & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) |
      (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_2_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_4_0[4]))));
  assign nor_539_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[4])
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1);
  assign nor_540_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1!=2'b00));
  assign MAC_1_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_51_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_51_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_51_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_1_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_36_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_36_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_36_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_2_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_3_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_36_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_2_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_3_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_50_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_96_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_50_nl);
  assign operator_ac_float_cctor_m_36_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_96_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_2_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_29_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_101_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_29_nl);
  assign operator_ac_float_cctor_m_36_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_101_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_2_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_2_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6[4]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_3_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6[4])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_51_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_2_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_3_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_38_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_74_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_38_nl);
  assign operator_ac_float_cctor_m_51_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_74_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_2_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_24_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_92_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_24_nl);
  assign operator_ac_float_cctor_m_51_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_92_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_2_ssc);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      | nor_540_cse);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
      | nor_539_cse);
  assign nor_541_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1!=2'b00));
  assign or_865_ssc = nor_541_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0;
  assign operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_4 = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1[0])
      & or_865_ssc;
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_2_nl = ~ or_865_ssc;
  assign operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_3_0 = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2,
      4'b1111, ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_2_nl);
  assign nor_542_cse = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]!=2'b00));
  assign or_866_nl = nor_542_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0;
  assign operator_ac_float_cctor_e_21_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[4:0]),
      or_866_nl);
  assign MAC_1_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_21_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_21_lpi_1_dfm_1_5_0!=6'b000000));
  assign MAC_1_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_6_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_6_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6[4]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6[4])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_36_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_36_nl);
  assign operator_ac_float_cctor_m_6_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_31_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_31_nl);
  assign operator_ac_float_cctor_m_6_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_ssc);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1 =
      conv_s2s_11_12({(~ operator_ac_float_cctor_m_21_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_21_lpi_1_dfm_1_5_0)})
      + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_2_ssc = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_3_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
      | nor_542_cse);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
      | nor_541_cse);
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_14_lpi_1_dfm) - $signed(operator_ac_float_cctor_e_29_lpi_1_dfm);
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_19_lpi_1_dfm) - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0);
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0
      = (z_out_3[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0[1:0];
  assign nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1[5:4]) + 2'b01;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0
      = nl_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0[1:0];
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0
      = (z_out_2[5:4]) + 2'b01;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0
      = nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0[1:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_15_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_14_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_13_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_12_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_47_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_47_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_47_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_46_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_47_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_17_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_17_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6[4])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_37_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_37_nl);
  assign operator_ac_float_cctor_m_17_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_33_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_33_nl);
  assign operator_ac_float_cctor_m_17_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_ssc);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_11_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_46_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_46_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_46_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_42_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_43_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0[4])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_16_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_16_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_ssc = (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6[4])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_44_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_44_nl);
  assign operator_ac_float_cctor_m_16_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_32_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_32_nl);
  assign operator_ac_float_cctor_m_16_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_ssc);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_10_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp = ~((operator_ac_float_cctor_m_60_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_60_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_60_lpi_1_dfm_1_3_0!=4'b0000));
  assign MAC_10_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp = ~((operator_ac_float_cctor_m_45_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_45_lpi_1_dfm_1_5_0!=6'b000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_38_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_39_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0[4])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_38_ssc = (~
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0[4]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_39_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0[4])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_10_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_10_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign or_887_nl = and_dcpl_1547 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm);
  assign operator_ac_float_cctor_e_15_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
      or_887_nl);
  assign or_889_nl = and_dcpl_1557 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm);
  assign operator_ac_float_cctor_e_30_lpi_1_dfm_mx0 = MUX_v_5_2_2(5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
      or_889_nl);
  assign MAC_10_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp = ~((operator_ac_float_cctor_m_30_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_30_lpi_1_dfm_1_5_0!=6'b000000));
  assign MAC_10_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp = ~((operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6!=5'b00000)
      | (operator_ac_float_cctor_m_15_lpi_1_dfm_1_5_4!=2'b00) | (operator_ac_float_cctor_m_15_lpi_1_dfm_1_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_ssc = (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_ssc = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0[4])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1
      = conv_s2s_11_12({(~ operator_ac_float_cctor_m_30_lpi_1_dfm_1_10_6) , (~ operator_ac_float_cctor_m_30_lpi_1_dfm_1_5_0)})
      + 12'b000000000001;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1 = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[11:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_38_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_39_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0[4])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_10_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1_5_0[5:4]!=2'b00))));
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_14_lpi_1_dfm) - $signed(operator_ac_float_cctor_e_33_lpi_1_dfm);
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_31_lpi_1_dfm) - $signed(operator_ac_float_cctor_e_63_lpi_1_dfm);
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_19_lpi_1_dfm) - $signed(operator_ac_float_cctor_e_34_lpi_1_dfm);
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2)
      - $signed(operator_ac_float_cctor_e_64_lpi_1_dfm);
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0)
      - $signed(operator_ac_float_cctor_e_65_lpi_1_dfm);
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp
      = $signed(operator_ac_float_cctor_e_29_lpi_1_dfm) - $signed(operator_ac_float_cctor_e_3_lpi_1_dfm);
  assign nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2) + 7'b0000001;
  assign MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1) + 7'b0000001;
  assign MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_16 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_17 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5:4]==2'b01));
  assign nl_MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0)
      + 7'b0000001;
  assign MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0)
      + 7'b0000001;
  assign MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0)
      + 7'b0000001;
  assign MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1)
      + 7'b0000001;
  assign MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0)
      + 7'b0000001;
  assign MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1) + 7'b0000001;
  assign MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]))})
      + conv_u2s_4_7(MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1) + 7'b0000001;
  assign MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2) + 7'b0000001;
  assign MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1) + 7'b0000001;
  assign MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1) + 7'b0000001;
  assign MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0)
      + 7'b0000001;
  assign MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0)
      + 7'b0000001;
  assign MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0)
      + 7'b0000001;
  assign MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign operator_i_e_1_lpi_1_dfm_mx0 = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[4:0]),
      5'b01111, and_dcpl_1579);
  assign nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl
      =  -conv_s2s_5_6(operator_i_e_1_lpi_1_dfm_mx0);
  assign MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl =
      nl_MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl[5:0];
  assign MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1
      = readslicef_6_1_5(MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl);
  assign nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl
      =  -conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse);
  assign MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl =
      nl_MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl[5:0];
  assign MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1
      = readslicef_6_1_5(MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_18 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]==2'b01));
  assign nl_MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0)
      + 7'b0000001;
  assign MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0)
      + 7'b0000001;
  assign MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1) + 7'b0000001;
  assign MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2) + 7'b0000001;
  assign MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0)
      + 7'b0000001;
  assign MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1) + 7'b0000001;
  assign MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0)
      + 7'b0000001;
  assign MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0)
      + 7'b0000001;
  assign MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6
      = readslicef_7_1_6(MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0)
      + 7'b0000001;
  assign MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_19 = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_22 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_28 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_26 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_32 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_36 = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_38 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_40 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_42 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5:4]==2'b01));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_48_mx0 = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0, MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0)})
      + 6'b000001;
  assign MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      nl_MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_49_mx0 = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0, MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva);
  assign MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_61_lpi_1_dfm);
  assign MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva);
  assign MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_62_lpi_1_dfm);
  assign nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0)})
      + 6'b000001;
  assign MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      nl_MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_63_lpi_1_dfm);
  assign MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva);
  assign MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_64_lpi_1_dfm);
  assign nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0)})
      + 6'b000001;
  assign MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      nl_MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_65_lpi_1_dfm);
  assign MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva);
  assign MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_14_lpi_1_dfm);
  assign MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva);
  assign MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp =
      $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_19_lpi_1_dfm);
  assign nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0)})
      + 6'b000001;
  assign MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_29_lpi_1_dfm);
  assign nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0)
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1)}) + 6'b000001;
  assign MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_3_lpi_1_dfm);
  assign nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0)
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1)}) + 6'b000001;
  assign MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_31_lpi_1_dfm);
  assign MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0);
  assign MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2);
  assign nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      + conv_s2s_5_6({(~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4)
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0)}) + 6'b000001;
  assign MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_33_lpi_1_dfm);
  assign MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva);
  assign MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(operator_i_e_1_lpi_1_dfm_mx0) - $signed(operator_ac_float_cctor_e_34_lpi_1_dfm);
  assign MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = $signed(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva);
  assign nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = conv_s2s_5_6(operator_i_e_1_lpi_1_dfm_mx0) + conv_s2s_5_6({(~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0)
      , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1)})
      + 6'b000001;
  assign MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp
      = nl_MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16 = ~((i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6[5:4]==2'b01));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16 = ~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6[5:4]==2'b01));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_4 =
      MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4[0]),
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_4, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_3_0
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0,
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_4 =
      MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4[0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_3_0
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_4 =
      MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4[0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_3_0
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4[1]);
  assign nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl
      = nl_MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl[6:0];
  assign MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1
      = readslicef_7_1_6(MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl);
  assign nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0
      + conv_s2s_5_6({1'b1 , (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0)})
      + 6'b000001;
  assign MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm =
      nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm[5:0];
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp = MUX_v_6_2_2(6'b110000,
      MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm, MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl
      = ({1'b1 , (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]))})
      + conv_u2s_4_7(MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)
      + 7'b0000001;
  assign MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl
      = nl_MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl[6:0];
  assign MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1
      = readslicef_7_1_6(MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_nl);
  assign nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1
      + conv_s2s_5_6({1'b1 , (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0)})
      + 6'b000001;
  assign MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl = nl_MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl[5:0];
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp = MUX_v_6_2_2(6'b110000,
      MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_nl, MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign and_dcpl_2 = ~((fsm_output[6:5]!=2'b00));
  assign or_tmp_20 = (fsm_output[1:0]!=2'b00);
  assign mux_tmp_31 = MUX_s_1_2_2((~ (fsm_output[1])), (fsm_output[1]), fsm_output[0]);
  assign nor_98_cse = ~((fsm_output[3:2]!=2'b00));
  assign mux_tmp_56 = MUX_s_1_2_2((~ (fsm_output[5])), (fsm_output[5]), fsm_output[4]);
  assign nor_tmp_6 = (fsm_output[5:4]==2'b11);
  assign not_tmp_212 = ~((fsm_output[5:4]!=2'b00));
  assign mux_tmp_65 = MUX_s_1_2_2(not_tmp_212, nor_tmp_6, fsm_output[1]);
  assign or_dcpl_193 = or_361_cse | (fsm_output[2]);
  assign or_dcpl_194 = (fsm_output[5]) | (fsm_output[1]);
  assign or_dcpl_195 = (fsm_output[6]) | (fsm_output[4]);
  assign or_dcpl_196 = or_dcpl_195 | or_dcpl_194;
  assign or_dcpl_197 = or_dcpl_196 | or_dcpl_193;
  assign and_dcpl_164 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_166 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_167 = (fsm_output[6]) & (~ (fsm_output[4]));
  assign and_dcpl_169 = and_dcpl_167 & (~ (fsm_output[5])) & and_dcpl_166;
  assign or_dcpl_200 = (~ (fsm_output[0])) | (fsm_output[3]);
  assign or_dcpl_201 = or_dcpl_200 | (~ (fsm_output[2]));
  assign or_dcpl_204 = (~ (fsm_output[6])) | (fsm_output[4]) | or_dcpl_194 | or_dcpl_201;
  assign and_dcpl_182 = nor_469_cse & (~ (fsm_output[2]));
  assign and_dcpl_183 = ~((fsm_output[5]) | (fsm_output[1]));
  assign and_dcpl_184 = ~((fsm_output[6]) | (fsm_output[4]));
  assign and_dcpl_185 = and_dcpl_184 & and_dcpl_183;
  assign and_dcpl_186 = and_dcpl_185 & and_dcpl_182;
  assign and_dcpl_187 = (~ (fsm_output[5])) & (fsm_output[1]);
  assign and_dcpl_188 = and_dcpl_184 & and_dcpl_187;
  assign and_dcpl_189 = and_dcpl_188 & and_dcpl_182;
  assign or_dcpl_207 = or_dcpl_195 | (fsm_output[5]);
  assign and_dcpl_190 = (fsm_output[0]) & (~ (fsm_output[3]));
  assign and_dcpl_191 = and_dcpl_190 & (fsm_output[2]);
  assign and_dcpl_192 = and_dcpl_185 & and_dcpl_191;
  assign and_dcpl_193 = nor_469_cse & (fsm_output[2]);
  assign and_dcpl_194 = and_dcpl_188 & and_dcpl_193;
  assign and_dcpl_195 = and_dcpl_188 & and_dcpl_191;
  assign and_dcpl_196 = (~ (fsm_output[0])) & (fsm_output[3]);
  assign and_dcpl_197 = and_dcpl_196 & (~ (fsm_output[2]));
  assign and_dcpl_198 = and_dcpl_185 & and_dcpl_197;
  assign and_dcpl_199 = and_dcpl_185 & and_dcpl_193;
  assign and_dcpl_200 = ~((fsm_output[5]) | (fsm_output[3]));
  assign xor_dcpl = (fsm_output[1]) ^ (fsm_output[0]);
  assign and_dcpl_202 = and_dcpl_184 & xor_dcpl;
  assign and_dcpl_203 = and_dcpl_202 & and_dcpl_200 & (fsm_output[2]);
  assign and_dcpl_206 = and_dcpl_184 & (~ (fsm_output[5]));
  assign and_dcpl_208 = and_dcpl_190 & (~ (fsm_output[2]));
  assign and_dcpl_209 = and_dcpl_188 & and_dcpl_208;
  assign and_dcpl_210 = (fsm_output[0]) & (fsm_output[3]);
  assign and_dcpl_211 = and_dcpl_210 & (~ (fsm_output[2]));
  assign and_dcpl_212 = and_dcpl_185 & and_dcpl_211;
  assign or_tmp_98 = (~((fsm_output[5:3]!=3'b000))) | (fsm_output[6]);
  assign or_tmp_100 = not_tmp_212 | (fsm_output[6]);
  assign mux_tmp_98 = MUX_s_1_2_2((~ (fsm_output[6])), (fsm_output[6]), or_6_cse);
  assign mux_tmp_99 = MUX_s_1_2_2(mux_tmp_98, or_tmp_100, fsm_output[3]);
  assign mux_106_nl = MUX_s_1_2_2(mux_tmp_99, or_tmp_98, fsm_output[2]);
  assign and_dcpl_213 = (~ mux_106_nl) & and_dcpl_166;
  assign or_tmp_102 = (fsm_output[0]) | (fsm_output[1]) | (fsm_output[6]);
  assign mux_tmp_101 = MUX_s_1_2_2(mux_tmp_98, or_dcpl_207, fsm_output[1]);
  assign or_tmp_104 = (fsm_output[1:0]!=2'b00) | mux_tmp_98;
  assign mux_113_nl = MUX_s_1_2_2(mux_8_cse, or_tmp_98, fsm_output[2]);
  assign and_dcpl_215 = (~ mux_113_nl) & and_1628_cse;
  assign and_dcpl_218 = and_dcpl_184 & and_dcpl_200 & ((~ (fsm_output[0])) | (fsm_output[2]))
      & (fsm_output[1]);
  assign or_tmp_107 = (~ (fsm_output[1])) | (fsm_output[5]) | (fsm_output[4]) | (fsm_output[6]);
  assign nand_nl = ~((fsm_output[1]) & (~ mux_tmp_98));
  assign mux_117_nl = MUX_s_1_2_2(nand_nl, or_tmp_107, fsm_output[0]);
  assign mux_118_nl = MUX_s_1_2_2(mux_117_nl, or_467_cse, fsm_output[3]);
  assign mux_114_nl = MUX_s_1_2_2(or_dcpl_207, or_tmp_100, fsm_output[1]);
  assign mux_115_nl = MUX_s_1_2_2(mux_114_nl, or_dcpl_196, fsm_output[0]);
  assign mux_116_nl = MUX_s_1_2_2(mux_115_nl, or_467_cse, fsm_output[3]);
  assign mux_119_itm = MUX_s_1_2_2(mux_118_nl, mux_116_nl, fsm_output[2]);
  assign or_319_nl = (fsm_output[0]) | mux_tmp_101;
  assign mux_122_nl = MUX_s_1_2_2(or_319_nl, or_tmp_102, fsm_output[3]);
  assign mux_120_nl = MUX_s_1_2_2(mux_tmp_98, or_dcpl_207, or_tmp_20);
  assign mux_121_nl = MUX_s_1_2_2(mux_120_nl, or_tmp_102, fsm_output[3]);
  assign mux_123_itm = MUX_s_1_2_2(mux_122_nl, mux_121_nl, fsm_output[2]);
  assign and_dcpl_220 = not_tmp_212 & (~ (fsm_output[3]));
  assign mux_102_nl = MUX_s_1_2_2(and_1628_cse, (~ or_tmp_20), fsm_output[2]);
  assign and_dcpl_222 = mux_102_nl & (~ (fsm_output[6])) & and_dcpl_220;
  assign and_dcpl_223 = and_dcpl_167 & and_dcpl_183;
  assign or_tmp_111 = (fsm_output[1]) | mux_tmp_98;
  assign or_323_nl = (fsm_output[1:0]!=2'b00) | or_tmp_100;
  assign mux_tmp_121 = MUX_s_1_2_2(or_tmp_104, or_323_nl, fsm_output[3]);
  assign and_dcpl_227 = and_dcpl_185 & and_dcpl_208;
  assign mux_145_nl = MUX_s_1_2_2(or_tmp_20, (fsm_output[3]), fsm_output[2]);
  assign and_dcpl_231 = (~ mux_145_nl) & and_dcpl_206;
  assign mux_146_nl = MUX_s_1_2_2(xor_dcpl, or_tmp_20, fsm_output[3]);
  assign mux_147_nl = MUX_s_1_2_2(mux_146_nl, (fsm_output[3]), fsm_output[2]);
  assign and_dcpl_232 = (~ mux_147_nl) & and_dcpl_206;
  assign mux_tmp_143 = MUX_s_1_2_2(nor_137_cse, (fsm_output[1]), fsm_output[2]);
  assign and_dcpl_243 = and_dcpl_202 & and_dcpl_200 & (~ (fsm_output[2]));
  assign mux_tmp_146 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[5]);
  assign mux_tmp_147 = MUX_s_1_2_2(not_tmp_212, mux_tmp_146, fsm_output[1]);
  assign and_245_nl = (fsm_output[1]) & mux_tmp_146;
  assign mux_154_nl = MUX_s_1_2_2(and_245_nl, mux_tmp_147, fsm_output[0]);
  assign mux_tmp_149 = MUX_s_1_2_2(mux_154_nl, nor_tmp_6, fsm_output[3]);
  assign mux_tmp_150 = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_tmp_20);
  assign not_tmp_284 = ~(and_1628_cse | (fsm_output[5:4]!=2'b00));
  assign or_51_nl = (fsm_output[3]) | (~ and_1628_cse);
  assign mux_161_nl = MUX_s_1_2_2(or_tmp_20, or_51_nl, fsm_output[2]);
  assign and_dcpl_245 = (~ mux_161_nl) & and_dcpl_206;
  assign and_dcpl_248 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_251 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_254 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_257 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign or_tmp_131 = (fsm_output[1:0]!=2'b10);
  assign mux_175_nl = MUX_s_1_2_2((~ or_tmp_131), or_tmp_20, fsm_output[2]);
  assign and_dcpl_260 = mux_175_nl & (~ (fsm_output[6])) & and_dcpl_220;
  assign mux_182_nl = MUX_s_1_2_2(or_dcpl_196, mux_tmp_101, fsm_output[0]);
  assign or_8_nl = (fsm_output[1]) | (fsm_output[6]);
  assign mux_181_nl = MUX_s_1_2_2(or_dcpl_196, or_8_nl, fsm_output[0]);
  assign mux_183_nl = MUX_s_1_2_2(mux_182_nl, mux_181_nl, fsm_output[3]);
  assign mux_178_nl = MUX_s_1_2_2(or_tmp_100, or_dcpl_207, fsm_output[1]);
  assign mux_179_nl = MUX_s_1_2_2(or_tmp_107, mux_178_nl, fsm_output[0]);
  assign or_57_nl = (fsm_output[1]) | (~ (fsm_output[0])) | (fsm_output[6]);
  assign mux_180_nl = MUX_s_1_2_2(mux_179_nl, or_57_nl, fsm_output[3]);
  assign mux_184_itm = MUX_s_1_2_2(mux_183_nl, mux_180_nl, fsm_output[2]);
  assign and_dcpl_277 = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_280 = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (~ (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]));
  assign and_dcpl_281 = and_dcpl_210 & (fsm_output[2]);
  assign and_dcpl_282 = and_dcpl_185 & and_dcpl_281;
  assign and_dcpl_283 = (~ (fsm_output[6])) & (fsm_output[4]);
  assign and_dcpl_284 = and_dcpl_283 & and_dcpl_183;
  assign and_dcpl_285 = and_dcpl_284 & and_dcpl_208;
  assign and_dcpl_286 = and_dcpl_284 & and_dcpl_191;
  assign and_dcpl_287 = and_dcpl_284 & and_dcpl_211;
  assign and_dcpl_288 = and_dcpl_284 & and_dcpl_281;
  assign and_dcpl_289 = (fsm_output[5]) & (~ (fsm_output[1]));
  assign and_dcpl_290 = and_dcpl_184 & and_dcpl_289;
  assign and_dcpl_291 = and_dcpl_290 & and_dcpl_208;
  assign and_dcpl_292 = and_dcpl_290 & and_dcpl_191;
  assign and_dcpl_293 = and_dcpl_290 & and_dcpl_211;
  assign and_dcpl_294 = and_dcpl_290 & and_dcpl_281;
  assign and_dcpl_295 = and_dcpl_283 & and_dcpl_289;
  assign and_dcpl_296 = and_dcpl_295 & and_dcpl_208;
  assign and_dcpl_297 = and_dcpl_295 & and_dcpl_191;
  assign and_dcpl_298 = and_dcpl_295 & and_dcpl_211;
  assign and_dcpl_299 = and_dcpl_295 & and_dcpl_281;
  assign and_dcpl_300 = and_dcpl_223 & and_dcpl_208;
  assign and_dcpl_327 = and_dcpl_185 & (~ (fsm_output[0])) & (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_345 = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign mux_tmp_188 = MUX_s_1_2_2(nor_tmp_6, (fsm_output[5]), fsm_output[1]);
  assign not_tmp_307 = ~((fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]));
  assign mux_tmp_223 = MUX_s_1_2_2((~ and_1628_cse), (fsm_output[1]), fsm_output[3]);
  assign or_dcpl_229 = or_dcpl_196 | or_dcpl_200 | (fsm_output[2]);
  assign and_dcpl_361 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_364 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_367 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_370 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_373 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_376 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_379 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_382 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_385 = and_dcpl_185 & (~ (fsm_output[0])) & (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_388 = and_dcpl_185 & (~((fsm_output[0]) | (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign and_dcpl_392 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_395 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_399 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_402 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_405 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_408 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_409 = and_dcpl_183 & and_dcpl_164;
  assign nor_177_nl = ~((~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[0]));
  assign or_386_nl = (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[0]);
  assign mux_tmp_236 = MUX_s_1_2_2(nor_177_nl, or_386_nl, MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_420 = and_dcpl_185 & and_dcpl_190 & (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[2]);
  assign and_dcpl_423 = and_dcpl_185 & and_dcpl_190 & (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & (fsm_output[2]);
  assign and_dcpl_426 = and_dcpl_185 & (~ (fsm_output[0])) & (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_429 = and_dcpl_185 & (~((fsm_output[0]) | (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign and_dcpl_432 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_dcpl_435 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign and_dcpl_452 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_455 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign or_tmp_153 = nor_137_cse | (fsm_output[4]);
  assign or_tmp_154 = (fsm_output[1]) | (~ (fsm_output[4]));
  assign and_dcpl_478 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_481 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign and_dcpl_482 = (fsm_output[0]) & (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_484 = and_dcpl_185 & and_dcpl_482 & and_dcpl_164;
  assign and_dcpl_485 = (fsm_output[0]) & (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]));
  assign and_dcpl_487 = and_dcpl_185 & and_dcpl_485 & and_dcpl_164;
  assign and_dcpl_496 = and_dcpl_188 & (fsm_output[0]) & (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign and_dcpl_499 = and_dcpl_188 & (fsm_output[0]) & (~ (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & nor_98_cse;
  assign and_dcpl_521 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_524 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign nor_tmp_26 = (fsm_output[1]) & (fsm_output[4]);
  assign mux_tmp_247 = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[1]);
  assign and_dcpl_552 = and_dcpl_185 & (fsm_output[0]) & (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_555 = and_dcpl_185 & (fsm_output[0]) & (~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_164;
  assign mux_261_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, and_2663_cse);
  assign mux_260_nl = MUX_s_1_2_2(mux_tmp_146, mux_tmp_188, fsm_output[3]);
  assign mux_262_nl = MUX_s_1_2_2(mux_261_nl, mux_260_nl, fsm_output[2]);
  assign and_dcpl_574 = ~(mux_262_nl | (fsm_output[6]));
  assign mux_tmp_257 = MUX_s_1_2_2((~ (fsm_output[4])), nor_tmp_26, fsm_output[3]);
  assign and_dcpl_596 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_599 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign mux_tmp_261 = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, fsm_output[1]);
  assign mux_268_nl = MUX_s_1_2_2(mux_tmp_147, mux_tmp_261, fsm_output[3]);
  assign mux_266_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, fsm_output[3]);
  assign mux_269_nl = MUX_s_1_2_2(mux_268_nl, mux_266_nl, fsm_output[2]);
  assign and_dcpl_624 = ~(mux_269_nl | (fsm_output[6]));
  assign and_dcpl_633 = (~ (fsm_output[0])) & (fsm_output[2]);
  assign nor_tmp_29 = (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[1]);
  assign and_dcpl_637 = and_dcpl_2 & (fsm_output[2]);
  assign and_dcpl_640 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_647 = and_dcpl_283 & and_dcpl_187;
  assign and_dcpl_654 = (fsm_output[5]) & (fsm_output[1]);
  assign and_dcpl_655 = and_dcpl_184 & and_dcpl_654;
  assign and_dcpl_663 = (fsm_output[3:2]==2'b11);
  assign and_dcpl_669 = and_dcpl_283 & and_dcpl_654;
  assign and_dcpl_679 = and_dcpl_167 & and_dcpl_187;
  assign and_dcpl_689 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_692 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign and_dcpl_720 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_723 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign and_dcpl_799 = and_dcpl_185 & (fsm_output[0]) & (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_802 = and_dcpl_185 & (fsm_output[0]) & (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_164;
  assign and_dcpl_854 = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign and_dcpl_857 = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign and_dcpl_937 = and_dcpl_206 & (~ or_tmp_131);
  assign and_dcpl_963 = and_dcpl_166 & and_dcpl_640;
  assign and_dcpl_964 = and_dcpl_206 & or_966_cse;
  assign and_dcpl_976 = and_dcpl_187 & (fsm_output[0]) & nor_98_cse;
  assign and_dcpl_981 = and_1628_cse & (~ (fsm_output[3]));
  assign and_dcpl_985 = nor_137_cse & and_dcpl_640;
  assign and_dcpl_990 = and_dcpl_206 & nor_137_cse;
  assign or_dcpl_257 = or_tmp_107 | or_dcpl_193;
  assign or_tmp_238 = ac_float_cctor_operator_return_63_sva | (~ and_dcpl_482);
  assign and_dcpl_1012 = and_dcpl_183 & (fsm_output[0]) & and_dcpl_164;
  assign or_dcpl_262 = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5:4]!=2'b01);
  assign and_dcpl_1017 = and_dcpl_206 & and_1628_cse;
  assign mux_362_nl = MUX_s_1_2_2(mux_tmp_99, mux_8_cse, fsm_output[2]);
  assign and_dcpl_1036 = (~ mux_362_nl) & nor_137_cse;
  assign and_dcpl_1054 = and_dcpl_183 & (~ (fsm_output[0])) & and_dcpl_164;
  assign and_dcpl_1070 = and_dcpl_206 & or_967_cse;
  assign and_dcpl_1077 = and_dcpl_187 & (~ (fsm_output[0]));
  assign and_dcpl_1078 = and_dcpl_1077 & and_dcpl_663;
  assign and_dcpl_1082 = and_dcpl_1077 & nor_98_cse;
  assign and_dcpl_1090 = and_dcpl_1077 & and_dcpl_640;
  assign and_dcpl_1097 = and_dcpl_654 & (~ (fsm_output[0]));
  assign and_dcpl_1098 = and_dcpl_1097 & nor_98_cse;
  assign and_dcpl_1102 = and_dcpl_1097 & and_dcpl_164;
  assign and_dcpl_1106 = and_dcpl_1097 & and_dcpl_640;
  assign and_dcpl_1110 = and_dcpl_1097 & and_dcpl_663;
  assign and_dcpl_1138 = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]!=2'b01));
  assign and_dcpl_1142 = and_dcpl_206 & and_dcpl_166;
  assign and_dcpl_1173 = and_dcpl_206 & or_968_cse;
  assign and_dcpl_1187 = and_dcpl_206 & ((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]!=2'b01));
  assign and_dcpl_1218 = and_dcpl_206 & (fsm_output[2:1]==2'b10);
  assign mux_385_nl = MUX_s_1_2_2(nor_tmp_6, mux_tmp_146, fsm_output[1]);
  assign mux_tmp_380 = MUX_s_1_2_2(mux_385_nl, mux_tmp_188, fsm_output[3]);
  assign and_dcpl_1267 = and_dcpl_640 & ((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0!=2'b01));
  assign nor_8_nl = ~((fsm_output[3]) | (~ (fsm_output[1])));
  assign mux_tmp_384 = MUX_s_1_2_2(nor_tmp_6, mux_tmp_146, nor_8_nl);
  assign mux_81_nl = MUX_s_1_2_2(mux_tmp_65, and_1593_cse, fsm_output[0]);
  assign mux_398_nl = MUX_s_1_2_2(not_tmp_307, mux_81_nl, fsm_output[3]);
  assign mux_tmp_393 = MUX_s_1_2_2(mux_398_nl, mux_80_cse, fsm_output[2]);
  assign nor_195_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[5:4]!=2'b00));
  assign or_tmp_275 = nor_195_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm)
      | (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]);
  assign or_608_nl = (~ (fsm_output[3])) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00);
  assign mux_tmp_402 = MUX_s_1_2_2(or_608_nl, or_tmp_275, fsm_output[2]);
  assign and_dcpl_1355 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[5:4]!=2'b00));
  assign or_tmp_291 = (~ (fsm_output[3])) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b01);
  assign and_dcpl_1363 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1366 = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]!=2'b01));
  assign and_dcpl_1369 = and_dcpl_206 & (fsm_output[0]) & (~ (fsm_output[2]));
  assign and_dcpl_1374 = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]!=2'b01));
  assign nor_199_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5:4]!=2'b00));
  assign or_tmp_300 = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
      | (fsm_output[3]) | nor_199_cse | (fsm_output[1:0]!=2'b00);
  assign nor_200_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp[5:4]!=2'b00));
  assign or_tmp_303 = nor_200_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp[6])
      | (~(MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs &
      (fsm_output[1:0]==2'b11)));
  assign and_dcpl_1383 = and_dcpl_640 & or_dcpl_262;
  assign and_dcpl_1389 = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5:4]!=2'b01));
  assign and_dcpl_1395 = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]!=2'b01));
  assign and_dcpl_1398 = and_dcpl_184 & (~((fsm_output[5]) | (fsm_output[2])));
  assign nor_203_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp[5:4]!=2'b00));
  assign or_tmp_319 = nor_203_cse | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp[6])
      | (~ and_1628_cse);
  assign not_tmp_606 = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp[5:4]!=2'b00))
      & (fsm_output[1:0]==2'b11));
  assign and_dcpl_1413 = and_dcpl_640 & or_730_cse;
  assign and_dcpl_1425 = and_dcpl_188 & and_dcpl_197;
  assign and_dcpl_1426 = and_dcpl_196 & (fsm_output[2]);
  assign and_dcpl_1427 = and_dcpl_188 & and_dcpl_1426;
  assign and_dcpl_1428 = and_dcpl_647 & and_dcpl_182;
  assign and_dcpl_1429 = and_dcpl_647 & and_dcpl_193;
  assign and_dcpl_1430 = and_dcpl_647 & and_dcpl_197;
  assign and_dcpl_1431 = and_dcpl_647 & and_dcpl_1426;
  assign and_dcpl_1432 = and_dcpl_655 & and_dcpl_182;
  assign and_dcpl_1433 = and_dcpl_655 & and_dcpl_193;
  assign and_dcpl_1434 = and_dcpl_655 & and_dcpl_197;
  assign and_dcpl_1435 = and_dcpl_655 & and_dcpl_1426;
  assign and_dcpl_1436 = and_dcpl_669 & and_dcpl_182;
  assign and_dcpl_1437 = and_dcpl_669 & and_dcpl_193;
  assign and_dcpl_1438 = and_dcpl_669 & and_dcpl_197;
  assign and_dcpl_1439 = and_dcpl_669 & and_dcpl_1426;
  assign and_dcpl_1440 = and_dcpl_679 & and_dcpl_182;
  assign and_dcpl_1450 = and_dcpl_206 & (~(or_tmp_131 | (fsm_output[3])));
  assign and_dcpl_1463 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5:4]!=2'b00));
  assign or_760_nl = ac_float_cctor_operator_return_59_sva | (~ (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | (fsm_output[1]);
  assign mux_tmp_477 = MUX_s_1_2_2(or_760_nl, (fsm_output[1]), MAC_11_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp);
  assign mux_tmp_481 = MUX_s_1_2_2((~ nor_tmp_26), or_900_cse, fsm_output[0]);
  assign or_763_nl = (fsm_output[0]) | (~ nor_tmp_26);
  assign mux_488_nl = MUX_s_1_2_2(or_763_nl, mux_tmp_481, nor_75_cse);
  assign mux_tmp_483 = MUX_s_1_2_2(mux_488_nl, mux_tmp_481, ac_float_cctor_operator_return_30_sva);
  assign and_dcpl_1547 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1550 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1551 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1554 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1557 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1562 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1565 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1568 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5:4]!=2'b00));
  assign and_dcpl_1575 = and_dcpl_185 & (~ (fsm_output[0])) & (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_dcpl_1578 = and_dcpl_185 & (~((fsm_output[0]) | (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign or_dcpl_485 = or_361_cse | (~ (fsm_output[2]));
  assign or_dcpl_486 = or_dcpl_196 | or_dcpl_485;
  assign or_dcpl_507 = or_dcpl_196 | or_dcpl_201;
  assign or_dcpl_509 = or_tmp_107 | or_dcpl_485;
  assign and_dcpl_1579 = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]==2'b01);
  assign return_imag_e_rsci_idat_mx0c1 = and_dcpl_169 & and_dcpl_164 & (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp[5:4]==2'b01)
      & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign return_real_e_rsci_idat_mx0c1 = and_dcpl_169 & and_dcpl_164 & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp[5:4]==2'b01);
  assign mux_157_nl = MUX_s_1_2_2(not_tmp_284, mux_tmp_150, fsm_output[3]);
  assign mux_158_nl = MUX_s_1_2_2(mux_157_nl, mux_tmp_149, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_mx0c2
      = ~(mux_158_nl | (fsm_output[6]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c1
      = and_dcpl_188 & nor_469_cse & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c2
      = and_dcpl_188 & nor_469_cse & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c3
      = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c4
      = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1[1])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3
      = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4
      = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1[1])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6
      = and_dcpl_185 & (~((fsm_output[0]) | (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3
      = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4
      = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1[1])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6
      = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (~ (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]));
  assign mux_230_nl = MUX_s_1_2_2(or_1078_cse, (~ mux_tmp_223), fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1
      = mux_230_nl & and_dcpl_206;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
      = mux_tmp_236 & and_dcpl_184 & and_dcpl_409;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
      = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
      = and_dcpl_185 & and_dcpl_190 & (fsm_output[2]) & (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
      = and_dcpl_185 & nor_469_cse & (fsm_output[2]) & (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
      = (~ mux_tmp_236) & and_dcpl_184 & and_dcpl_409;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
      = and_dcpl_185 & and_dcpl_190 & (fsm_output[2]) & (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2])))
      & nor_98_cse;
  assign or_920_nl = (~ (fsm_output[3])) | (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[0]) | (~ and_1593_cse);
  assign or_921_nl = (fsm_output[3]) | (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[5]) | (fsm_output[4]);
  assign mux_291_nl = MUX_s_1_2_2(or_920_nl, or_921_nl, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4
      = ~(mux_291_nl | (fsm_output[6]));
  assign nor_295_nl = ~((MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      | (~ (fsm_output[0])) | (fsm_output[1]) | (fsm_output[4]));
  assign nor_296_nl = ~((MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[0]) | (~ nor_tmp_26));
  assign mux_292_nl = MUX_s_1_2_2(nor_295_nl, nor_296_nl, fsm_output[3]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5
      = mux_292_nl & and_dcpl_637;
  assign or_922_nl = (~ (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[2]) | (~ (fsm_output[6]));
  assign or_923_nl = (~ (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_924_nl = (~ (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_303_nl = MUX_s_1_2_2(or_923_nl, or_924_nl, fsm_output[2]);
  assign mux_304_nl = MUX_s_1_2_2(or_922_nl, mux_303_nl, fsm_output[3]);
  assign or_925_nl = (~ (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_926_nl = (~ (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_301_nl = MUX_s_1_2_2(or_925_nl, or_926_nl, fsm_output[2]);
  assign or_927_nl = (~ (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_928_nl = (~ (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_300_nl = MUX_s_1_2_2(or_927_nl, or_928_nl, fsm_output[2]);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_300_nl, fsm_output[3]);
  assign mux_305_nl = MUX_s_1_2_2(mux_304_nl, mux_302_nl, fsm_output[5]);
  assign or_929_nl = (~ (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_930_nl = (~ (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_297_nl = MUX_s_1_2_2(or_929_nl, or_930_nl, fsm_output[2]);
  assign or_931_nl = (~ (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_932_nl = (~ (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_296_nl = MUX_s_1_2_2(or_931_nl, or_932_nl, fsm_output[2]);
  assign mux_298_nl = MUX_s_1_2_2(mux_297_nl, mux_296_nl, fsm_output[3]);
  assign or_933_nl = (~ (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_934_nl = (~ (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_294_nl = MUX_s_1_2_2(or_933_nl, or_934_nl, fsm_output[2]);
  assign or_935_nl = (~ (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_936_nl = (~ (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_293_nl = MUX_s_1_2_2(or_935_nl, or_936_nl, fsm_output[2]);
  assign mux_295_nl = MUX_s_1_2_2(mux_294_nl, mux_293_nl, fsm_output[3]);
  assign mux_299_nl = MUX_s_1_2_2(mux_298_nl, mux_295_nl, fsm_output[5]);
  assign mux_306_nl = MUX_s_1_2_2(mux_305_nl, mux_299_nl, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8
      = ~(mux_306_nl | or_tmp_131);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9
      = and_dcpl_188 & (~((fsm_output[0]) | (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10
      = and_dcpl_188 & (~((fsm_output[0]) | (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21
      = and_dcpl_679 & (~((fsm_output[0]) | (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2])))
      & nor_98_cse;
  assign or_937_nl = (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[6]));
  assign or_938_nl = (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_325_nl = MUX_s_1_2_2(or_937_nl, or_938_nl, fsm_output[3]);
  assign or_939_nl = (~ (fsm_output[3])) | (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_326_nl = MUX_s_1_2_2(mux_325_nl, or_939_nl, fsm_output[2]);
  assign or_940_nl = (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_941_nl = (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_323_nl = MUX_s_1_2_2(or_940_nl, or_941_nl, fsm_output[3]);
  assign or_942_nl = (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_943_nl = (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_322_nl = MUX_s_1_2_2(or_942_nl, or_943_nl, fsm_output[3]);
  assign mux_324_nl = MUX_s_1_2_2(mux_323_nl, mux_322_nl, fsm_output[2]);
  assign mux_327_nl = MUX_s_1_2_2(mux_326_nl, mux_324_nl, fsm_output[5]);
  assign or_944_nl = (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_945_nl = (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_319_nl = MUX_s_1_2_2(or_944_nl, or_945_nl, fsm_output[3]);
  assign or_946_nl = (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_947_nl = (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_318_nl = MUX_s_1_2_2(or_946_nl, or_947_nl, fsm_output[3]);
  assign mux_320_nl = MUX_s_1_2_2(mux_319_nl, mux_318_nl, fsm_output[2]);
  assign or_948_nl = (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_949_nl = (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_316_nl = MUX_s_1_2_2(or_948_nl, or_949_nl, fsm_output[3]);
  assign or_950_nl = (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign or_951_nl = (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[6]);
  assign mux_315_nl = MUX_s_1_2_2(or_950_nl, or_951_nl, fsm_output[3]);
  assign mux_317_nl = MUX_s_1_2_2(mux_316_nl, mux_315_nl, fsm_output[2]);
  assign mux_321_nl = MUX_s_1_2_2(mux_320_nl, mux_317_nl, fsm_output[5]);
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, mux_321_nl, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7
      = ~(mux_328_nl | or_tmp_131);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8
      = and_dcpl_188 & (~ (fsm_output[0])) & (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9
      = and_dcpl_647 & (~ (fsm_output[0])) & (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10
      = and_dcpl_647 & (~ (fsm_output[0])) & (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11
      = and_dcpl_647 & (~ (fsm_output[0])) & (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12
      = and_dcpl_647 & and_dcpl_196 & (fsm_output[2]) & (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13
      = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14
      = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15
      = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16
      = and_dcpl_655 & (~ (fsm_output[0])) & (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17
      = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18
      = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19
      = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20
      = and_dcpl_669 & (~ (fsm_output[0])) & (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21
      = and_dcpl_679 & (~ (fsm_output[0])) & (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2])))
      & nor_98_cse;
  assign nand_46_nl = ~((MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[6]));
  assign or_952_nl = (~ (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_346_nl = MUX_s_1_2_2(nand_46_nl, or_952_nl, fsm_output[3]);
  assign or_953_nl = (~ (fsm_output[3])) | (~ (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_347_nl = MUX_s_1_2_2(mux_346_nl, or_953_nl, fsm_output[2]);
  assign or_954_nl = (~ (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_955_nl = (~ (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_344_nl = MUX_s_1_2_2(or_954_nl, or_955_nl, fsm_output[3]);
  assign or_956_nl = (~ (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_957_nl = (~ (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_343_nl = MUX_s_1_2_2(or_956_nl, or_957_nl, fsm_output[3]);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, mux_343_nl, fsm_output[2]);
  assign mux_348_nl = MUX_s_1_2_2(mux_347_nl, mux_345_nl, fsm_output[5]);
  assign or_958_nl = (~ (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_959_nl = (~ (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_340_nl = MUX_s_1_2_2(or_958_nl, or_959_nl, fsm_output[3]);
  assign or_960_nl = (~ (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_961_nl = (~ (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_339_nl = MUX_s_1_2_2(or_960_nl, or_961_nl, fsm_output[3]);
  assign mux_341_nl = MUX_s_1_2_2(mux_340_nl, mux_339_nl, fsm_output[2]);
  assign or_962_nl = (~ (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_963_nl = (~ (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_337_nl = MUX_s_1_2_2(or_962_nl, or_963_nl, fsm_output[3]);
  assign or_964_nl = (~ (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign or_965_nl = (~ (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[6]);
  assign mux_336_nl = MUX_s_1_2_2(or_964_nl, or_965_nl, fsm_output[3]);
  assign mux_338_nl = MUX_s_1_2_2(mux_337_nl, mux_336_nl, fsm_output[2]);
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, mux_338_nl, fsm_output[5]);
  assign mux_349_nl = MUX_s_1_2_2(mux_348_nl, mux_342_nl, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8
      = ~(mux_349_nl | or_tmp_131);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9
      = and_dcpl_188 & (~((fsm_output[0]) | (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10
      = and_dcpl_188 & (~((fsm_output[0]) | (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13
      = and_dcpl_647 & (~((fsm_output[0]) | (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14
      = and_dcpl_647 & and_dcpl_196 & (fsm_output[2]) & (~ (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18
      = and_dcpl_655 & (~((fsm_output[0]) | (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22
      = and_dcpl_669 & (~((fsm_output[0]) | (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_663;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23
      = and_dcpl_679 & (~((fsm_output[0]) | (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0
      = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2])
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1
      = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2])))
      & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c1
      = (((MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_1_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_1_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_1_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_1_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c3
      = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5:4]!=2'b01))
      & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c4
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c3
      = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5:4]!=2'b01))
      & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c4
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c1
      = (((~ MAC_4_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) &
      (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_4_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c2
      = and_dcpl_206 & (MAC_4_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp
      | (~ (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])))
      & and_dcpl_981 & (~((fsm_output[2]) | MAC_4_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign mux_358_nl = MUX_s_1_2_2(and_dcpl_485, (fsm_output[0]), ac_float_cctor_operator_return_63_sva);
  assign mux_359_nl = MUX_s_1_2_2(mux_358_nl, or_tmp_238, MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign nor_389_nl = ~(ac_float_cctor_operator_return_48_sva | (~ mux_359_nl));
  assign mux_357_nl = MUX_s_1_2_2(or_tmp_238, (~ (fsm_output[0])), ac_float_cctor_operator_return_48_sva);
  assign mux_360_nl = MUX_s_1_2_2(nor_389_nl, mux_357_nl, ac_float_cctor_operator_return_42_sva);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c3
      = mux_360_nl & and_dcpl_206 & (~ or_1078_cse) & (fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c4
      = and_dcpl_206 & ((~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_48_sva) & nor_137_cse & (~ ac_float_cctor_operator_return_42_sva)
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c5
      = (((MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_63_sva)) | ac_float_cctor_operator_return_48_sva)
      & and_dcpl_184 & and_dcpl_1012;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c6
      = and_dcpl_1017 & and_dcpl_164 & or_dcpl_262;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c7
      = and_dcpl_1017 & and_dcpl_164 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5:4]==2'b01);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c3
      = and_dcpl_1017 & and_dcpl_164 & or_730_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c4
      = and_dcpl_1017 & and_dcpl_164 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[5:4]==2'b01);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c1
      = (((MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_3_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_3_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_3_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_3_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c3
      = (((~ ac_float_cctor_operator_return_60_sva) & (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_12_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_1054;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c4
      = and_dcpl_206 & (ac_float_cctor_operator_return_60_sva | (~ (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])))
      & nor_137_cse & (fsm_output[3:2]==2'b01) & (~ MAC_12_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c5
      = (((MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_62_sva)) | ac_float_cctor_operator_return_42_sva)
      & and_dcpl_184 & and_dcpl_1012;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c6
      = and_dcpl_206 & ((~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_62_sva) & and_dcpl_166 & (~ ac_float_cctor_operator_return_42_sva)
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c7
      = and_dcpl_1070 & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c8
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign nor_393_nl = ~((MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[6])));
  assign mux_374_nl = MUX_s_1_2_2(nor_393_nl, (fsm_output[6]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm);
  assign nor_395_nl = ~((fsm_output[2]) | (~ mux_374_nl));
  assign nor_396_nl = ~((~((~ (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)) | (fsm_output[6]));
  assign nor_397_nl = ~((~(MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      | (~ (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_373_nl = MUX_s_1_2_2(nor_396_nl, nor_397_nl, fsm_output[2]);
  assign mux_375_nl = MUX_s_1_2_2(nor_395_nl, mux_373_nl, fsm_output[3]);
  assign nor_398_nl = ~((~(MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_399_nl = ~((~(MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      | (~ (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_371_nl = MUX_s_1_2_2(nor_398_nl, nor_399_nl, fsm_output[2]);
  assign nor_400_nl = ~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm
      | (~ (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_401_nl = ~((~(MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_370_nl = MUX_s_1_2_2(nor_400_nl, nor_401_nl, fsm_output[2]);
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, mux_370_nl, fsm_output[3]);
  assign mux_376_nl = MUX_s_1_2_2(mux_375_nl, mux_372_nl, fsm_output[5]);
  assign nor_402_nl = ~((~(MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_403_nl = ~((~(MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_367_nl = MUX_s_1_2_2(nor_402_nl, nor_403_nl, fsm_output[2]);
  assign nor_404_nl = ~((~(MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_405_nl = ~((~((~ (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)) | (fsm_output[6]));
  assign mux_366_nl = MUX_s_1_2_2(nor_404_nl, nor_405_nl, fsm_output[2]);
  assign mux_368_nl = MUX_s_1_2_2(mux_367_nl, mux_366_nl, fsm_output[3]);
  assign nor_406_nl = ~((~(MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      | (~ (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_407_nl = ~((~(MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_364_nl = MUX_s_1_2_2(nor_406_nl, nor_407_nl, fsm_output[2]);
  assign nor_408_nl = ~((~(MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      | (~ (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign nor_409_nl = ~((~(MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      | (~ (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[6]));
  assign mux_363_nl = MUX_s_1_2_2(nor_408_nl, nor_409_nl, fsm_output[2]);
  assign mux_365_nl = MUX_s_1_2_2(mux_364_nl, mux_363_nl, fsm_output[3]);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, mux_365_nl, fsm_output[5]);
  assign mux_377_nl = MUX_s_1_2_2(mux_376_nl, mux_369_nl, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c9
      = mux_377_nl & (~(or_tmp_131 | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c10
      = (((MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1078;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c11
      = (((MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1082;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c12
      = (((MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1077 & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c13
      = (((MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1090;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c14
      = (((MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)) |
      MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1078;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c15
      = (((MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1098;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c16
      = (((MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)) |
      MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1102;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c17
      = (((MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1106;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c18
      = (((MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1110;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c19
      = (((MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1098;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c20
      = (((MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1102;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c21
      = (((MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1106;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c22
      = (((MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_283 & and_dcpl_1110;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c23
      = (((MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm))
      | MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp)
      & and_dcpl_167 & and_dcpl_1082;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c5
      = and_dcpl_1138 & and_dcpl_963;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c6
      = and_dcpl_1142 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c1
      = (((MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_5_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_5_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_5_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_1628_cse
      & (~ MAC_5_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & nor_98_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c3
      = and_dcpl_990 & (((~ MAC_10_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)
      & (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_10_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c4
      = and_dcpl_990 & and_dcpl_164 & (~ MAC_10_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp)
      & (MAC_10_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp | (~
      (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c5
      = (((MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_3_sva)) | ac_float_cctor_operator_return_29_sva)
      & and_dcpl_184 & and_dcpl_1012;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c6
      = and_dcpl_206 & ((~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_3_sva) & and_dcpl_166 & (~ ac_float_cctor_operator_return_29_sva)
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c7
      = and_dcpl_1173 & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c8
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c5
      = and_dcpl_1187 & and_dcpl_963;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c6
      = and_dcpl_1142 & (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c1
      = (((MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_6_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_6_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_6_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_6_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c3
      = (((MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_29_sva)) | MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp)
      & and_dcpl_184 & and_dcpl_1054;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c4
      = and_dcpl_206 & ((~ (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_29_sva) & nor_137_cse & (~ MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp)
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c5
      = and_dcpl_1218 & (((~ ac_float_cctor_operator_return_31_sva) & (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_12_sva) & and_dcpl_190;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c6
      = and_dcpl_1218 & and_dcpl_190 & (~ ac_float_cctor_operator_return_12_sva)
      & (ac_float_cctor_operator_return_31_sva | (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c7
      = and_dcpl_964 & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c8
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c1
      = (((MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_7_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_7_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_7_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_7_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c3
      = (((~ ac_float_cctor_operator_return_30_sva) & (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp) & and_dcpl_184
      & and_dcpl_1054;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c4
      = and_dcpl_206 & (ac_float_cctor_operator_return_30_sva | (~ (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & nor_137_cse & (~ MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp)
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c5
      = (((~ ac_float_cctor_operator_return_32_sva) & (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_17_sva) & and_dcpl_184 & and_dcpl_1012;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c6
      = and_dcpl_206 & (ac_float_cctor_operator_return_32_sva | (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & (~((fsm_output[3]) | (~ (fsm_output[0])) | (fsm_output[1]))) & (~ ac_float_cctor_operator_return_17_sva)
      & (fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c7
      = and_dcpl_990 & and_dcpl_1267;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c8
      = and_dcpl_990 & and_dcpl_640 & (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0==2'b01);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0
      = and_dcpl_188 & nor_469_cse & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1
      = and_dcpl_188 & nor_469_cse & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c1
      = (((MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & (~ MAC_8_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp)) |
      MAC_8_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_184
      & and_dcpl_976;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c2
      = and_dcpl_206 & ((~ (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      | MAC_8_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp) & and_dcpl_981
      & (~((fsm_output[2]) | MAC_8_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c3
      = and_dcpl_1218 & (((~ ac_float_cctor_operator_return_17_sva) & (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | ac_float_cctor_operator_return_12_sva) & nor_469_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c4
      = and_dcpl_1218 & nor_469_cse & (~ ac_float_cctor_operator_return_12_sva) &
      (ac_float_cctor_operator_return_17_sva | (~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c5
      = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5:4]!=2'b01))
      & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c6
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
      = and_dcpl_188 & nor_469_cse & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
      = and_dcpl_188 & nor_469_cse & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c3
      = and_dcpl_206 & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5:4]!=2'b01))
      & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c4
      = and_dcpl_990 & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5:4]==2'b01)
      & and_dcpl_640;
  assign or_610_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00);
  assign mux_409_nl = MUX_s_1_2_2((~ and_1628_cse), or_610_nl, fsm_output[3]);
  assign mux_410_nl = MUX_s_1_2_2(mux_409_nl, or_tmp_275, fsm_output[2]);
  assign or_609_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[5:4]!=2'b00);
  assign mux_411_nl = MUX_s_1_2_2(mux_tmp_402, mux_410_nl, or_609_nl);
  assign or_605_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6]);
  assign mux_412_nl = MUX_s_1_2_2(mux_411_nl, mux_tmp_402, or_605_nl);
  assign operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c1 = (~ mux_412_nl) & and_dcpl_206;
  assign operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm))
      & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c3 = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
      | nor_195_cse) & and_dcpl_184 & and_dcpl_1054;
  assign operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c4 = and_dcpl_1138 & and_dcpl_985;
  assign nor_429_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp[5:4]!=2'b00));
  assign nor_431_nl = ~(nor_429_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp[6])
      | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm
      & (fsm_output[1:0]==2'b11))));
  assign nor_432_nl = ~((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00));
  assign mux_413_nl = MUX_s_1_2_2(nor_431_nl, nor_432_nl, fsm_output[3]);
  assign nor_433_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
      | and_dcpl_1355 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (fsm_output[3]) | (fsm_output[0]) | (fsm_output[1]));
  assign mux_414_nl = MUX_s_1_2_2(mux_413_nl, nor_433_nl, fsm_output[2]);
  assign operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c1 = mux_414_nl & and_dcpl_206;
  assign operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c2 = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_16_tmp[6])
      | nor_429_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c3 = (and_dcpl_1355 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0)
      & and_dcpl_184 & and_dcpl_1054;
  assign operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c4 = and_dcpl_1187 & and_dcpl_985;
  assign or_633_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b01);
  assign mux_415_nl = MUX_s_1_2_2((~ and_1628_cse), or_633_nl, fsm_output[3]);
  assign or_632_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp[5:4]!=2'b00);
  assign mux_416_nl = MUX_s_1_2_2(or_tmp_291, mux_415_nl, or_632_nl);
  assign or_630_nl = (~ ac_float_cctor_operator_return_17_sva) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp[6]);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, or_tmp_291, or_630_nl);
  assign or_629_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm)
      | (fsm_output[3]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      | and_dcpl_1363 | (fsm_output[1:0]!=2'b00);
  assign mux_418_nl = MUX_s_1_2_2(mux_417_nl, or_629_nl, fsm_output[2]);
  assign operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c1 = (~ mux_418_nl) & and_dcpl_206;
  assign operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_16_tmp[6])
      | (~ ac_float_cctor_operator_return_17_sva)) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c3 = (and_dcpl_1363 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm))
      & and_dcpl_184 & and_dcpl_1054;
  assign operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c4 = and_dcpl_1366 & and_dcpl_963;
  assign nor_438_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp[6])
      | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp[5:4]!=2'b00))
      & (fsm_output[1]))));
  assign nor_439_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1]));
  assign mux_419_nl = MUX_s_1_2_2(nor_438_nl, nor_439_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c1 = mux_419_nl & and_dcpl_1369;
  assign operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_30_tmp[6]))
      & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c3 = and_dcpl_1374 & and_dcpl_963;
  assign nor_56_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[5:4]!=2'b01));
  assign or_652_nl = (fsm_output[3]) | or_tmp_303;
  assign mux_422_nl = MUX_s_1_2_2(or_652_nl, or_tmp_300, fsm_output[2]);
  assign or_354_nl = (fsm_output[1:0]!=2'b01);
  assign mux_420_nl = MUX_s_1_2_2(or_tmp_303, or_354_nl, fsm_output[3]);
  assign mux_421_nl = MUX_s_1_2_2(mux_420_nl, or_tmp_300, fsm_output[2]);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, mux_421_nl, nor_56_cse);
  assign operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c1 = (~ mux_423_nl) & and_dcpl_206;
  assign operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c2 = ((~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_20_tmp[6])
      | nor_200_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c3 = (nor_199_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm))
      & and_dcpl_184 & and_dcpl_1054;
  assign operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c4 = and_dcpl_1142 & and_dcpl_1383;
  assign nor_442_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp[5:4]!=2'b00));
  assign nor_443_nl = ~(nor_442_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp[6])
      | (~(MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs &
      (fsm_output[1]))));
  assign nor_444_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1]));
  assign mux_424_nl = MUX_s_1_2_2(nor_443_nl, nor_444_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c1 = mux_424_nl & and_dcpl_1369;
  assign operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c2 = ((~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_24_tmp[6])
      | nor_442_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c3 = and_dcpl_1389 & and_dcpl_963;
  assign nor_447_nl = ~((~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp[6])
      | (~(((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp[5:4]!=2'b00))
      & (fsm_output[1]))));
  assign nor_448_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1]));
  assign mux_425_nl = MUX_s_1_2_2(nor_447_nl, nor_448_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c1 = mux_425_nl & and_dcpl_1369;
  assign operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp[5:4]!=2'b00)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_26_tmp[6])
      | (~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c3 = and_dcpl_1395 & and_dcpl_963;
  assign nor_450_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp[5:4]!=2'b00));
  assign nor_451_nl = ~(nor_450_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp[6])
      | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm
      & (fsm_output[1:0]==2'b11))));
  assign nor_452_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00));
  assign mux_426_nl = MUX_s_1_2_2(nor_451_nl, nor_452_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c1 = mux_426_nl & and_dcpl_1398;
  assign operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c2 = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_20_tmp[6])
      | nor_450_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c3 = and_dcpl_1374 & and_dcpl_985;
  assign or_680_nl = (fsm_output[3]) | or_tmp_319;
  assign mux_427_nl = MUX_s_1_2_2(or_tmp_319, or_tmp_20, fsm_output[3]);
  assign mux_428_nl = MUX_s_1_2_2(or_680_nl, mux_427_nl, nor_56_cse);
  assign operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c1 = (~ mux_428_nl) & and_dcpl_1398;
  assign operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c2 = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_22_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm)
      | nor_203_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c3 = and_dcpl_990 & and_dcpl_1383;
  assign or_687_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp[6])
      | not_tmp_606;
  assign mux_429_nl = MUX_s_1_2_2(or_687_nl, or_tmp_20, fsm_output[3]);
  assign or_686_nl = (fsm_output[3]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp[6])
      | not_tmp_606;
  assign mux_430_nl = MUX_s_1_2_2(mux_429_nl, or_686_nl, or_730_cse);
  assign operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c1 = (~ mux_430_nl) & and_dcpl_1398;
  assign operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_24_tmp[6]))
      & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c3 = and_dcpl_990 & and_dcpl_1413;
  assign nor_456_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp[5:4]!=2'b00));
  assign nor_457_nl = ~(nor_456_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp[6])
      | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm
      & (fsm_output[1:0]==2'b11))));
  assign nor_458_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00));
  assign mux_431_nl = MUX_s_1_2_2(nor_457_nl, nor_458_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c1 = mux_431_nl & and_dcpl_1398;
  assign operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c2 = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_26_tmp[6])
      | nor_456_cse) & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c3 = and_dcpl_1389 & and_dcpl_985;
  assign nor_461_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp[6])
      | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp[5:4]!=2'b00))
      & (fsm_output[1:0]==2'b11))));
  assign nor_462_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]!=2'b01)
      | (fsm_output[1:0]!=2'b00));
  assign mux_432_nl = MUX_s_1_2_2(nor_461_nl, nor_462_nl, fsm_output[3]);
  assign operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c1 = mux_432_nl & and_dcpl_1398;
  assign operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c2 = ((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp[5:4]!=2'b00)))
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_28_tmp[6]))
      & and_dcpl_184 & and_dcpl_976;
  assign operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c3 = and_dcpl_1395 & and_dcpl_985;
  assign or_dcpl_526 = (and_dcpl_195 & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_6_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_198 & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_14_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_527 = (and_dcpl_195 & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_198 & (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_528 = (and_dcpl_198 & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_15_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_195 & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_7_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_529 = (and_dcpl_198 & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_195 & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_530 = (and_dcpl_195 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_8_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_198 & MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_16_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_531 = (and_dcpl_195 & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_198 & (~ MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_532 = (and_dcpl_195 & MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_2_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_198 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_11_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_533 = (and_dcpl_195 & (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | (and_dcpl_198 & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_534 = (and_dcpl_198 & MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_12_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_195 & MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_3_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_535 = (and_dcpl_198 & (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | (and_dcpl_195 & (~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs));
  assign or_dcpl_536 = (and_dcpl_195 & MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_4_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6))
      | (and_dcpl_198 & MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_13_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6));
  assign or_dcpl_537 = (and_dcpl_195 & (~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_198 & (~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs));
  assign or_dcpl_538 = (and_dcpl_198 & MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_10_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (and_dcpl_195 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_9_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign or_dcpl_539 = (and_dcpl_198 & (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_195 & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_540 = (and_dcpl_198 & MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_14_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (and_dcpl_195 & MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_5_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign or_dcpl_541 = (and_dcpl_198 & (~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_195 & (~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs));
  assign or_dcpl_543 = (((and_dcpl_195 & (~ MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (and_dcpl_194 & (~ MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)))
      & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) |
      (and_dcpl_198 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_10_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign mux_nl = MUX_s_1_2_2(and_dcpl_195, and_dcpl_212, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign or_1030_nl = (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | and_dcpl_212;
  assign mux_517_nl = MUX_s_1_2_2(mux_nl, or_1030_nl, and_dcpl_194);
  assign or_dcpl_544 = mux_517_nl | (and_dcpl_198 & (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs));
  assign nor_567_nl = ~(MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      | (~ and_dcpl_212));
  assign nor_568_nl = ~(MAC_3_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (~ and_dcpl_195));
  assign mux_518_nl = MUX_s_1_2_2(nor_567_nl, nor_568_nl, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign or_dcpl_546 = mux_518_nl | (and_dcpl_198 & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & (~ MAC_11_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs & and_dcpl_194
      & (~ MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign mux_519_nl = MUX_s_1_2_2(and_dcpl_195, and_dcpl_212, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign or_dcpl_548 = mux_519_nl | (and_dcpl_198 & (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | ((~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)
      & and_dcpl_194);
  assign or_dcpl_550 = (((and_dcpl_198 & (~ MAC_12_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (and_dcpl_194 & (~ MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)))
      & MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs) | (and_dcpl_195
      & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs & (~
      MAC_4_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign or_dcpl_551 = and_dcpl_198 | and_dcpl_194;
  assign or_dcpl_552 = (or_dcpl_551 & (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs))
      | (and_dcpl_195 & (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs));
  assign or_dcpl_554 = (((and_dcpl_198 & (~ MAC_13_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      | (and_dcpl_194 & (~ MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)))
      & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) |
      (and_dcpl_195 & MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
      & (~ MAC_5_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign or_dcpl_555 = (or_dcpl_551 & (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      | (and_dcpl_195 & (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs));
  assign or_dcpl_558 = ((MAC_1_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp
      | MAC_1_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp) & and_dcpl_209)
      | (and_dcpl_192 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs &
      and_dcpl_199);
  assign or_dcpl_577 = (and_dcpl_192 & MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)
      | (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs &
      and_dcpl_199);
  assign or_dcpl_578 = (and_dcpl_192 & MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs)
      | (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs &
      and_dcpl_199);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_ssc = and_dcpl_189
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_192 | and_dcpl_194 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c5
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c6;
  assign nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt
      = nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_2_cse = (~
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_3_cse = (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_4_cse = (~
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[5])) & and_dcpl_199;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_5_cse = (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[5])
      & and_dcpl_199;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_6_cse = (~
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_192;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_7_cse = (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_192;
  assign nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign and_1240_ssc = and_dcpl_1070 & and_dcpl_963;
  assign or_572_nl = (or_967_cse & (fsm_output[0])) | (fsm_output[1]);
  assign mux_387_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_572_nl);
  assign mux_388_nl = MUX_s_1_2_2(mux_tmp_261, mux_387_nl, fsm_output[3]);
  assign mux_389_nl = MUX_s_1_2_2(mux_388_nl, mux_tmp_380, fsm_output[2]);
  assign or_573_ssc = mux_389_nl | (fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_1_cse
      = (~ (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_192;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_2_cse
      = (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_192;
  assign nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt
      = nl_MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4:0];
  assign and_1282_ssc = and_dcpl_1173 & and_dcpl_963;
  assign or_581_nl = (or_968_cse & (fsm_output[0])) | (fsm_output[1]);
  assign mux_391_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_581_nl);
  assign mux_392_nl = MUX_s_1_2_2(mux_tmp_65, mux_391_nl, fsm_output[3]);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, mux_tmp_384, fsm_output[2]);
  assign or_582_ssc = mux_393_nl | (fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_6_cse
      = (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_192;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_7_cse
      = (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_192;
  assign and_dcpl_1740 = not_tmp_212 & nor_501_cse;
  assign and_1883_cse = and_dcpl_1740 & (fsm_output[2:0]==3'b010);
  assign and_1886_cse = and_dcpl_1740 & and_1628_cse & (~ (fsm_output[2]));
  assign and_1888_cse = and_dcpl_1740 & and_1628_cse & (fsm_output[2]);
  assign nor_578_cse = ~((fsm_output[2:0]!=3'b000));
  assign and_1893_cse = not_tmp_212 & (~ (fsm_output[6])) & (fsm_output[3]) & nor_578_cse;
  assign and_dcpl_1752 = (fsm_output[1:0]==2'b10);
  assign and_1899_cse = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2]));
  assign and_1909_cse = and_dcpl_1740 & and_dcpl_1752 & (fsm_output[2]);
  assign and_dcpl_1779 = not_tmp_212 & (~ (fsm_output[6])) & (fsm_output[3]);
  assign and_dcpl_1780 = and_dcpl_1779 & nor_578_cse;
  assign and_1925_cse = and_dcpl_1740 & (fsm_output[2:0]==3'b111);
  assign and_dcpl_1788 = and_dcpl_1779 & (fsm_output[2:0]==3'b001);
  assign and_dcpl_1857 = and_dcpl_1740 & and_dcpl_1752 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2])));
  assign and_dcpl_1860 = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2]);
  assign and_dcpl_1872 = and_dcpl_1740 & and_dcpl_1752 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2])));
  assign and_dcpl_1875 = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2]);
  assign and_dcpl_1885 = (fsm_output[3:0]==4'b0010);
  assign and_dcpl_1892 = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2])
      & (~ (fsm_output[4])) & and_dcpl_2 & and_dcpl_1885;
  assign and_dcpl_1939 = and_dcpl_1740 & and_dcpl_1752 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2])));
  assign and_dcpl_1942 = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2]);
  assign and_dcpl_1952 = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2])
      & (~ (fsm_output[4])) & and_dcpl_2 & and_dcpl_1885;
  assign and_dcpl_1962 = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2]);
  assign and_2125_cse = not_tmp_212 & nor_501_cse & (fsm_output[2:0]==3'b010);
  assign and_dcpl_1995 = and_dcpl_1740 & and_dcpl_1752 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2])));
  assign and_dcpl_1998 = and_dcpl_1740 & and_dcpl_1752 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2]);
  assign and_dcpl_2029 = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2])
      & (~ (fsm_output[4])) & and_dcpl_2 & and_dcpl_1885;
  assign and_2241_cse = not_tmp_212 & nor_501_cse & nor_137_cse & (fsm_output[2]);
  assign and_2261_cse = and_dcpl_1740 & nor_137_cse & (fsm_output[2]);
  assign and_2264_cse = and_dcpl_1740 & (fsm_output[2:0]==3'b101);
  assign and_2317_cse = not_tmp_212 & nor_501_cse & (fsm_output[2:0]==3'b101);
  assign and_2326_cse = not_tmp_212 & nor_501_cse & (fsm_output[2:0]==3'b110);
  assign and_2438_cse = not_tmp_212 & (~ (fsm_output[6])) & (fsm_output[3]) & (~
      (fsm_output[1])) & (fsm_output[0]) & (~ (fsm_output[2]));
  assign mux_526_nl = MUX_s_1_2_2(not_tmp_212, or_6_cse, fsm_output[6]);
  assign mux_527_nl = MUX_s_1_2_2(mux_526_nl, (fsm_output[6]), fsm_output[3]);
  assign mux_533_nl = MUX_s_1_2_2(or_tmp_100, (fsm_output[6]), fsm_output[3]);
  assign mux_528_nl = MUX_s_1_2_2(mux_527_nl, mux_533_nl, fsm_output[2]);
  assign and_dcpl_2475 = (~ mux_528_nl) & (fsm_output[1:0]==2'b11);
  assign nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_conc_32_itm_4_0 = MUX_v_5_2_2(MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
      MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      and_dcpl_199);
  assign nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl = MUX_v_5_2_2((MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_39_nl = ~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_39_nl);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_conc_29_itm_4_0 = MUX_v_5_2_2(MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl,
      and_dcpl_199);
  assign reg_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_1_cse
      = ~((and_dcpl_206 & and_dcpl_191) | and_dcpl_189);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse = (~
      and_dcpl_192) & (~((~(nor_137_cse ^ (fsm_output[2]))) | (fsm_output[6]))) &
      and_dcpl_220;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_5_cse = ~(and_dcpl_206
      & (fsm_output[3:1]==3'b011));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_90_cse = (~
      and_dcpl_194) & mux_tmp_143 & (~ (fsm_output[6])) & and_dcpl_220;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_71_cse = (~
      and_dcpl_199) & and_dcpl_222;
  assign mux_150_nl = MUX_s_1_2_2(or_tmp_20, and_1628_cse, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse = (~
      and_dcpl_199) & (~(mux_150_nl | (fsm_output[6]))) & and_dcpl_220;
  assign mux_151_nl = MUX_s_1_2_2(or_tmp_20, mux_tmp_31, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_cse = (~ and_dcpl_192)
      & (~(mux_151_nl | (fsm_output[6]))) & and_dcpl_220;
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0
      = conv_s2s_5_6(delay_lane_real_e_2_sva) + conv_s2s_5_6(taps_real_e_rsci_idat[19:15]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0
      = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0[5:0];
  assign or_735_nl = nor_478_cse | (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp[6])
      | (fsm_output[5:4]!=2'b00);
  assign mux_477_nl = MUX_s_1_2_2(or_6_cse, or_735_nl, and_1628_cse);
  assign or_733_nl = nor_479_cse | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
      | (fsm_output[5:4]!=2'b00);
  assign mux_475_nl = MUX_s_1_2_2(or_733_nl, or_6_cse, fsm_output[0]);
  assign mux_476_nl = MUX_s_1_2_2((~ mux_475_nl), mux_tmp_56, fsm_output[1]);
  assign mux_478_nl = MUX_s_1_2_2((~ mux_477_nl), mux_476_nl, fsm_output[2]);
  assign mux_472_nl = MUX_s_1_2_2(mux_tmp_56, nor_tmp_6, or_730_cse);
  assign mux_473_nl = MUX_s_1_2_2(mux_tmp_56, mux_472_nl, fsm_output[0]);
  assign or_729_nl = (fsm_output[2:1]!=2'b00);
  assign mux_474_nl = MUX_s_1_2_2(mux_473_nl, nor_tmp_6, or_729_nl);
  assign mux_479_nl = MUX_s_1_2_2(mux_478_nl, mux_474_nl, fsm_output[3]);
  assign or_736_rgt = mux_479_nl | (fsm_output[6]);
  assign and_1462_rgt = (nor_478_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_22_tmp[6])
      | (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
      & and_dcpl_184 & and_dcpl_976;
  assign and_1465_rgt = (nor_479_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm))
      & and_dcpl_184 & and_dcpl_1054;
  assign and_1466_rgt = and_dcpl_1142 & and_dcpl_1413;
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_14_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign and_1789_nl = and_dcpl_195 & nor_558_m1c;
  assign and_1790_nl = and_dcpl_198 & nor_558_m1c;
  assign mux1h_7_nl = MUX1HOT_v_6_4_2(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
      (z_out_21[5:0]), (z_out_7[5:0]), 6'b110000, {and_dcpl_186 , and_1789_nl , and_1790_nl
      , or_dcpl_540});
  assign not_1827_nl = ~ or_dcpl_541;
  assign and_1787_itm = MUX_v_6_2_2(6'b000000, mux1h_7_nl, not_1827_nl);
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0 = conv_s2s_5_6(delay_lane_imag_e_3_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[24:20]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0[5:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_33_cse = ~((~(and_dcpl_186 | and_dcpl_243
      | (~ mux_119_itm) | and_dcpl_194)) | and_dcpl_189);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0
      = conv_s2s_5_6(delay_lane_imag_e_2_sva) + conv_s2s_5_6(taps_imag_e_rsci_idat[19:15]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0[5:0];
  assign nor_474_tmp = ~((~(MAC_16_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp
      | (~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0
      = conv_s2s_5_6(delay_lane_real_e_2_sva) + conv_s2s_5_6(taps_imag_e_rsci_idat[19:15]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0[5:0];
  assign nor_495_tmp = ~((~((~ (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_3_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nor_774_cse = ~((fsm_output[2]) | (fsm_output[3]) | (fsm_output[5]));
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0
      = conv_s2s_5_6(delay_lane_imag_e_2_sva) + conv_s2s_5_6(taps_real_e_rsci_idat[19:15]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0[5:0];
  assign nor_493_tmp = ~((~(MAC_4_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp
      | (~ (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0
      = conv_s2s_5_6(delay_lane_imag_e_7_sva) + conv_s2s_5_6(taps_imag_e_rsci_idat[44:40]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0
      = nl_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0[5:0];
  assign nor_489_tmp = ~((~((~ (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_6_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0 = conv_s2s_5_6(delay_lane_real_e_7_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[44:40]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0[5:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_35_cse = ~((~(and_dcpl_186 | and_dcpl_243
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_194 | and_dcpl_215)) | and_dcpl_189);
  assign nor_487_tmp = ~((~((~ (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_7_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0 = conv_s2s_5_6(delay_lane_imag_e_7_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[44:40]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0[5:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_38_cse = operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_ssc
      & (~ and_dcpl_189);
  assign nor_485_tmp = ~((~((~ (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_8_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0 = conv_s2s_5_6(delay_lane_real_e_7_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[44:40]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0[5:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_41_cse = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_1_ssc
      & (~ and_dcpl_189);
  assign nor_519_tmp = ~((~((~ (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_1_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_1_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0 = conv_s2s_5_6(delay_lane_real_e_3_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[24:20]);
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0 = nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0[5:0];
  assign and_1785_m1c = and_dcpl_212 & nor_559_m1c;
  assign nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0 = conv_s2s_5_6(delay_lane_imag_e_4_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[29:25]);
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0 = nl_ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0[5:0];
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_ssc = and_dcpl_186 | and_dcpl_260
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_198;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse =
      and_dcpl_195 | and_dcpl_212;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse =
      and_dcpl_282 | and_dcpl_285;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse =
      and_dcpl_286 | and_dcpl_287;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse =
      and_dcpl_288 | and_dcpl_291;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse =
      and_dcpl_292 | and_dcpl_294;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse =
      and_dcpl_293 | and_dcpl_296;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse =
      and_dcpl_297 | and_dcpl_299;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse =
      and_dcpl_298 | and_dcpl_300;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0
      = conv_s2s_5_6(delay_lane_imag_e_5_sva) + conv_s2s_5_6(taps_imag_e_rsci_idat[34:30]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_1_ssc = and_dcpl_186
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4
      | and_dcpl_327 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6
      | and_dcpl_194 | and_dcpl_195 | and_dcpl_198 | and_dcpl_212;
  assign mux_561_cse = MUX_s_1_2_2((fsm_output[1]), (~ (fsm_output[1])), fsm_output[3]);
  assign nor_794_cse = ~((fsm_output[3]) | (~((fsm_output[1:0]!=2'b01))));
  assign nor_796_cse = ~((fsm_output[6:4]!=3'b000));
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0
      = conv_s2s_5_6(delay_lane_real_e_5_sva) + conv_s2s_5_6(taps_imag_e_rsci_idat[34:30]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_2_ssc = and_dcpl_186
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4
      | and_dcpl_345 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6
      | and_dcpl_194 | and_dcpl_195 | and_dcpl_198 | and_dcpl_212;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_26_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_2_ssc & (~ and_dcpl_574);
  assign nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = conv_s2s_5_6(delay_lane_imag_e_5_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[34:30]);
  assign MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_27_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_3_ssc & (~ and_dcpl_624);
  assign nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = conv_s2s_5_6(delay_lane_real_e_5_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[34:30]);
  assign MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = nl_MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:0];
  assign mux_289_nl = MUX_s_1_2_2(not_tmp_212, mux_tmp_261, fsm_output[3]);
  assign mux_288_nl = MUX_s_1_2_2(mux_tmp_147, nor_tmp_6, fsm_output[3]);
  assign mux_290_nl = MUX_s_1_2_2(mux_289_nl, mux_288_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_28_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_4_ssc & (mux_290_nl
      | (fsm_output[6]));
  assign nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm = conv_s2s_5_6(delay_lane_imag_e_6_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[39:35]);
  assign MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm = nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[5:0];
  assign mux_313_nl = MUX_s_1_2_2(not_tmp_212, nor_tmp_6, and_2663_cse);
  assign mux_312_nl = MUX_s_1_2_2(not_tmp_212, nor_tmp_6, fsm_output[3]);
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, mux_312_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_29_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_5_ssc & (mux_314_nl
      | (fsm_output[6]));
  assign nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = conv_s2s_5_6(delay_lane_real_e_6_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[39:35]);
  assign MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm = nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:0];
  assign mux_334_nl = MUX_s_1_2_2(not_tmp_212, and_1593_cse, fsm_output[3]);
  assign mux_335_nl = MUX_s_1_2_2(and_dcpl_220, mux_334_nl, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_30_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_6_ssc & (mux_335_nl
      | (fsm_output[6]));
  assign nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = conv_s2s_5_6(delay_lane_imag_e_6_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[39:35]);
  assign MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm = nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_31_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_7_ssc & (~((fsm_output[3])
      & (~ mux_tmp_143) & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_mx0c1));
  assign nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = conv_s2s_5_6(delay_lane_real_e_6_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[39:35]);
  assign MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm = nl_MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:0];
  assign mux_233_nl = MUX_s_1_2_2(xor_dcpl, or_tmp_20, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_44_cse = ~((~(((~(mux_233_nl | (fsm_output[6])))
      & and_dcpl_220) | and_dcpl_243 | and_dcpl_192)) | and_dcpl_189);
  assign nor_491_tmp = ~((~((~ (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_5_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) | MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_46_cse = operator_13_2_true_AC_TRN_AC_WRAP_1_or_5_ssc
      & (~ and_dcpl_189);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_48_cse = ~((~(and_dcpl_243 | and_dcpl_209
      | and_dcpl_192)) | and_dcpl_189);
  assign nor_476_tmp = ~((~(MAC_15_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp
      | (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_31_ssc = (~ nor_476_tmp) & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_32_ssc = nor_476_tmp & and_dcpl_209;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_2_ssc =
      and_dcpl_243 | and_dcpl_254 | and_dcpl_257 | and_dcpl_199 | and_dcpl_194 |
      and_dcpl_215;
  assign MAC_15_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1,
      MAC_15_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm
      = conv_s2s_6_7(MAC_15_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm =
      nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_3_ssc =
      and_dcpl_243 | and_dcpl_361 | and_dcpl_364 | and_dcpl_199 | and_dcpl_194 |
      and_dcpl_215;
  assign MAC_16_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1,
      MAC_16_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm
      = conv_s2s_6_7(MAC_16_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm =
      nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_4_ssc =
      and_dcpl_243 | and_dcpl_367 | and_dcpl_370 | and_dcpl_199 | and_dcpl_194;
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg)}) +
      7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_nl
      = ~((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_23_nl
      = ~(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_nl
      = MUX1HOT_v_7_3_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_acc_nl,
      7'b1110000, MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_nor_23_nl
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_itm
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_5_ssc =
      and_dcpl_243 | and_dcpl_373 | and_dcpl_376 | and_dcpl_199 | and_dcpl_194;
  assign MAC_10_r_ac_float_4_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4,
      MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign MAC_10_r_ac_float_4_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0,
      MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm
      = conv_s2s_6_7({MAC_10_r_ac_float_4_else_and_nl , MAC_10_r_ac_float_4_else_and_1_nl})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm =
      nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6:0];
  assign MAC_11_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0,
      MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt
      = conv_s2s_6_7(MAC_11_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt =
      nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_6_ssc =
      and_dcpl_243 | and_dcpl_379 | and_dcpl_382 | and_dcpl_385 | and_dcpl_388 |
      and_dcpl_192 | and_dcpl_195;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_7_ssc =
      and_dcpl_243 | and_dcpl_392 | and_dcpl_395 | and_dcpl_192 | and_dcpl_195;
  assign MAC_12_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1,
      MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm
      = conv_s2s_6_7(MAC_12_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm =
      nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc =
      and_dcpl_243 | and_dcpl_405 | and_dcpl_408 | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
      | and_dcpl_194;
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg)}) + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_15_sva_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_ssc
      = ~(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva[21]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      = ~((~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_nl
      = MUX1HOT_v_6_3_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5:0]),
      6'b110000, (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_ssc
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_itm
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_seb);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_ssc
      = and_dcpl_243 | and_dcpl_379 | and_dcpl_382 | and_dcpl_420 | and_dcpl_423
      | and_dcpl_194;
  assign MAC_10_r_ac_float_1_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4,
      MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign MAC_10_r_ac_float_1_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0,
      MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2s_6_7({MAC_10_r_ac_float_1_else_and_nl , MAC_10_r_ac_float_1_else_and_1_nl})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_ssc
      & (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_2_ssc
      = and_dcpl_243 | and_dcpl_392 | and_dcpl_395 | and_dcpl_426 | and_dcpl_429
      | and_dcpl_194;
  assign MAC_11_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0,
      MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2s_6_7(MAC_11_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_2_ssc
      & (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_3_ssc
      = and_dcpl_243 | and_dcpl_248 | and_dcpl_251 | and_dcpl_426 | and_dcpl_429
      | and_dcpl_192;
  assign MAC_12_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0,
      MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2s_6_7(MAC_12_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_3_ssc
      & (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_4_ssc
      = and_dcpl_243 | and_dcpl_432 | and_dcpl_435 | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
      | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
      | and_dcpl_194;
  assign MAC_13_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1,
      MAC_13_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2s_6_7(MAC_13_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_4_ssc
      & (~ and_dcpl_189);
  assign MAC_14_r_ac_float_1_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1,
      MAC_14_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt
      = conv_s2s_6_7(MAC_14_r_ac_float_1_else_and_nl) + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_5_ssc
      = and_dcpl_243 | and_dcpl_405 | and_dcpl_408 | and_dcpl_385 | and_dcpl_388
      | and_dcpl_194;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1
      | and_dcpl_720 | and_dcpl_723 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5
      | and_dcpl_195 | and_dcpl_198 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_1_ssc = and_dcpl_218 | and_dcpl_209
      | and_dcpl_199 | and_dcpl_198;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_6_ssc = and_dcpl_1450 | and_dcpl_209
      | and_dcpl_327 | and_dcpl_198;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_7_ssc = and_dcpl_1450 | and_dcpl_209
      | and_dcpl_345 | and_dcpl_198;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1
      = ~(and_2261_cse | and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_1_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1
      | and_dcpl_496 | and_dcpl_499;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_2_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1
      | and_dcpl_496 | and_dcpl_499;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_2_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1
      | and_dcpl_521 | and_dcpl_524 | and_dcpl_552 | and_dcpl_555 | and_dcpl_195;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_3_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_212;
  assign and_594_ssc = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2])
      & nor_98_cse;
  assign and_597_ssc = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2])))
      & nor_98_cse;
  assign and_606_ssc = and_dcpl_185 & (~ (fsm_output[0])) & (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_164;
  assign and_609_ssc = and_dcpl_185 & (~((fsm_output[0]) | (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])))
      & and_dcpl_164;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_5_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_212;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_6_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1
      | and_dcpl_209 | and_dcpl_212;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_1_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1
      | and_dcpl_720 | and_dcpl_723 | and_dcpl_799 | and_dcpl_802 | and_dcpl_198
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_7_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1
      | and_dcpl_209 | and_dcpl_199 | and_dcpl_212;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_2_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1
      | and_dcpl_478 | and_dcpl_481 | and_dcpl_799 | and_dcpl_802 | and_dcpl_195
      | and_dcpl_198 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_9_ssc = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
      | and_dcpl_209 | and_dcpl_212;
  assign and_537_ssc = and_dcpl_188 & (~ (fsm_output[0])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2])
      & nor_98_cse;
  assign and_540_ssc = and_dcpl_188 & (~((fsm_output[0]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2])))
      & nor_98_cse;
  assign and_543_ssc = and_dcpl_188 & and_dcpl_190 & (~ (fsm_output[2])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign and_546_ssc = and_dcpl_188 & and_dcpl_190 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1])));
  assign mux_459_nl = MUX_s_1_2_2((~ or_900_cse), nor_tmp_26, fsm_output[3]);
  assign nor_470_nl = ~(and_1628_cse | (fsm_output[4]));
  assign mux_458_nl = MUX_s_1_2_2(nor_470_nl, (fsm_output[4]), fsm_output[3]);
  assign mux_460_nl = MUX_s_1_2_2(mux_459_nl, mux_458_nl, fsm_output[2]);
  assign mux_254_nl = MUX_s_1_2_2(mux_tmp_247, nor_tmp_26, fsm_output[0]);
  assign mux_255_nl = MUX_s_1_2_2((~ (fsm_output[4])), mux_254_nl, fsm_output[3]);
  assign mux_252_nl = MUX_s_1_2_2((~ (fsm_output[4])), (fsm_output[4]), fsm_output[3]);
  assign mux_256_nl = MUX_s_1_2_2(mux_255_nl, mux_252_nl, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_ssc = (((~ mux_460_nl) & and_dcpl_2)
      | and_dcpl_192) & (~((~ mux_256_nl) & and_dcpl_2));
  assign operator_i_m_1_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_18});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl);
  assign operator_i_m_1_lpi_1_dfm_mx0w3_5_0 = MUX_v_6_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl,
      6'b111111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc);
  assign operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_54_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_55_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_54_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_55_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_54_nl);
  assign operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_54_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_55_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_106_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_nl);
  assign operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_106_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_54_ssc);
  assign operator_r_m_1_lpi_1_dfm_mx0w4_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_20});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_nl);
  assign operator_r_m_1_lpi_1_dfm_mx0w4_5_0 = MUX_v_6_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_nl,
      6'b111111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc);
  assign operator_i_m_8_lpi_1_dfm_mx0w10_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_28_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_44_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_22});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_71_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_44_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_71_nl);
  assign operator_i_m_8_lpi_1_dfm_mx0w10_5_4 = MUX_v_2_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl,
      2'b11, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_28_ssc);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_67_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_44_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_67_nl);
  assign operator_i_m_8_lpi_1_dfm_mx0w10_3_0 = MUX_v_4_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl,
      4'b1111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_28_ssc);
  assign operator_i_m_9_lpi_1_dfm_mx0w10_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_19});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_74_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_74_nl);
  assign operator_i_m_9_lpi_1_dfm_mx0w10_5_4 = MUX_v_2_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_56_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_68_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_68_nl);
  assign operator_i_m_9_lpi_1_dfm_mx0w10_3_0 = MUX_v_4_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_38);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_38);
  assign operator_r_m_4_lpi_1_dfm_mx0w5_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_38});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_91_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_54_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_91_nl);
  assign operator_r_m_4_lpi_1_dfm_mx0w5_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_54_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_80_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_80_nl);
  assign operator_r_m_4_lpi_1_dfm_mx0w5_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_62_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6[4])
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_36);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6[4])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_36);
  assign operator_r_m_14_lpi_1_dfm_mx0w5_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_36});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_84_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_84_nl);
  assign operator_r_m_14_lpi_1_dfm_mx0w5_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_63_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_81_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_81_nl);
  assign operator_r_m_14_lpi_1_dfm_mx0w5_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_55_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc);
  assign operator_r_m_6_lpi_1_dfm_mx0w5_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_5_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_11_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_32});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_93_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_11_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_49_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_93_nl);
  assign operator_r_m_6_lpi_1_dfm_mx0w5_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_49_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_5_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_75_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_11_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_67_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_75_nl);
  assign operator_r_m_6_lpi_1_dfm_mx0w5_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_67_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_5_ssc);
  assign operator_r_m_lpi_1_dfm_mx0w6_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_16});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_89_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_50_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_89_nl);
  assign operator_r_m_lpi_1_dfm_mx0w6_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_50_nl,
      2'b11, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_76_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_32_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_76_nl);
  assign operator_r_m_lpi_1_dfm_mx0w6_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_59_nl,
      4'b1111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_16_ssc);
  assign operator_r_m_2_lpi_1_dfm_mx0w6_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_42});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_88_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_51_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_88_nl);
  assign operator_r_m_2_lpi_1_dfm_mx0w6_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_51_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_77_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_36_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_77_nl);
  assign operator_r_m_2_lpi_1_dfm_mx0w6_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_20_ssc);
  assign operator_r_m_3_lpi_1_dfm_mx0w6_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_40});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_87_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_52_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_87_nl);
  assign operator_r_m_3_lpi_1_dfm_mx0w6_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_52_nl,
      2'b11, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_78_nl = ~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_38_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_78_nl);
  assign operator_r_m_3_lpi_1_dfm_mx0w6_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl,
      4'b1111, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_22_ssc);
  assign operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_62_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_63_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_52_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_64_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_52_nl);
  assign operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_64_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_62_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_16_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_104_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_16_nl);
  assign operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_104_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_62_ssc);
  assign operator_r_m_15_lpi_1_dfm_mx0w4_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_17});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_90_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_53_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_90_nl);
  assign operator_r_m_15_lpi_1_dfm_mx0w4_5_4 = MUX_v_2_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_53_nl,
      2'b11, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_79_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_34_ssc;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_79_nl);
  assign operator_r_m_15_lpi_1_dfm_mx0w4_3_0 = MUX_v_4_2_2(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl,
      4'b1111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_18_ssc);
  assign operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_50_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_51_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_55_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_51_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_65_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_55_nl);
  assign operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_65_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_50_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_17_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_51_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_107_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_17_nl);
  assign operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_107_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_50_ssc);
  assign operator_i_m_6_lpi_1_dfm_mx0w4_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_26});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_73_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_73_nl);
  assign operator_i_m_6_lpi_1_dfm_mx0w4_5_4 = MUX_v_2_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_57_nl,
      2'b11, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_69_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_40_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_69_nl);
  assign operator_i_m_6_lpi_1_dfm_mx0w4_3_0 = MUX_v_4_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_61_nl,
      4'b1111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_24_ssc);
  assign operator_i_m_7_lpi_1_dfm_mx0w3_10_6 = MUX1HOT_v_5_3_2(5'b01111, 5'b10000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0,
      {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_26_ssc
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_42_ssc , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_24});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_72_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_42_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_72_nl);
  assign operator_i_m_7_lpi_1_dfm_mx0w3_5_4 = MUX_v_2_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_58_nl,
      2'b11, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_26_ssc);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_70_nl = ~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_42_ssc;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_70_nl);
  assign operator_i_m_7_lpi_1_dfm_mx0w3_3_0 = MUX_v_4_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_60_nl,
      4'b1111, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_26_ssc);
  assign operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_58_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_59_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_53_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_59_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_66_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_53_nl);
  assign operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_66_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_58_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_18_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_59_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_105_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_18_nl);
  assign operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_105_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_58_ssc);
  assign operator_ac_float_cctor_m_1_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_62_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_63_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_33_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_33_nl);
  assign operator_ac_float_cctor_m_1_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_62_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_63_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_108_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_nl);
  assign operator_ac_float_cctor_m_1_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_108_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_62_ssc);
  assign operator_ac_float_cctor_m_35_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_58_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_59_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_16_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_59_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_64_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_16_nl);
  assign operator_ac_float_cctor_m_35_lpi_1_dfm_1_5_0 = MUX_v_6_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_64_nl,
      6'b111111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_58_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_30_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6[4]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_31_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6[4])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_43_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_30_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_31_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_48_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_72_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_48_nl);
  assign operator_ac_float_cctor_m_43_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_72_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_24_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_97_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_24_nl);
  assign operator_ac_float_cctor_m_43_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_97_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_8_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm);
  assign operator_ac_float_cctor_m_28_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_30_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_31_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_34_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_65_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_34_nl);
  assign operator_ac_float_cctor_m_28_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_65_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_17_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_31_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_109_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_17_nl);
  assign operator_ac_float_cctor_m_28_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_109_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_30_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_8_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1,
      ac_float_cctor_operator_return_12_sva);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_26_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6[4]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_27_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6[4])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_42_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_26_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_27_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_49_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_73_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_49_nl);
  assign operator_ac_float_cctor_m_42_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_73_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_25_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_98_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_25_nl);
  assign operator_ac_float_cctor_m_42_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_98_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm);
  assign operator_ac_float_cctor_m_27_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_26_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_27_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_35_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_66_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_35_nl);
  assign operator_ac_float_cctor_m_27_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_66_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_18_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_27_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_110_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_18_nl);
  assign operator_ac_float_cctor_m_27_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_110_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_26_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_7_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1,
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign operator_ac_float_cctor_m_41_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_22_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_23_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_44_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_67_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_44_nl);
  assign operator_ac_float_cctor_m_41_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_67_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_19_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_92_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_19_nl);
  assign operator_ac_float_cctor_m_41_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_92_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_6_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm);
  assign operator_ac_float_cctor_m_26_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_22_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_23_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_36_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_67_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_36_nl);
  assign operator_ac_float_cctor_m_26_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_67_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_19_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_23_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_111_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_19_nl);
  assign operator_ac_float_cctor_m_26_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_111_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_22_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_6_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1,
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign operator_ac_float_cctor_m_40_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_18_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_19_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_45_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_68_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_45_nl);
  assign operator_ac_float_cctor_m_40_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_68_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_20_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_93_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_20_nl);
  assign operator_ac_float_cctor_m_40_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_93_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_5_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_5_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1,
      ac_float_cctor_operator_return_63_sva);
  assign operator_ac_float_cctor_m_25_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_18_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_19_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_37_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_68_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_37_nl);
  assign operator_ac_float_cctor_m_25_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_68_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_20_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_19_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_112_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_20_nl);
  assign operator_ac_float_cctor_m_25_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_112_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_18_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_5_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1,
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_14_ssc = (~
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6[4]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_15_ssc = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6[4])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1;
  assign operator_ac_float_cctor_m_54_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6,
      5'b01111, 5'b10000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_15_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_25_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_75_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_25_nl);
  assign operator_ac_float_cctor_m_54_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_75_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_64_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_nl);
  assign operator_ac_float_cctor_m_54_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_64_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_4_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_4_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1,
      ac_float_cctor_operator_return_62_sva);
  assign operator_ac_float_cctor_m_24_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_38_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_69_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_38_nl);
  assign operator_ac_float_cctor_m_24_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_69_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_21_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_113_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_21_nl);
  assign operator_ac_float_cctor_m_24_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_113_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_4_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1,
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1,
      ac_float_cctor_operator_return_61_sva);
  assign operator_ac_float_cctor_m_23_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_10_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_11_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_28_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_70_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_28_nl);
  assign operator_ac_float_cctor_m_23_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_70_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_22_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_11_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_104_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_22_nl);
  assign operator_ac_float_cctor_m_23_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_104_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_10_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_3_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1,
      MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1,
      ac_float_cctor_operator_return_60_sva);
  assign operator_ac_float_cctor_m_22_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_6_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_7_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_29_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_71_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_29_nl);
  assign operator_ac_float_cctor_m_22_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_71_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_23_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_7_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_105_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_23_nl);
  assign operator_ac_float_cctor_m_22_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_105_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_6_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_2_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1,
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_4_0
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm);
  assign operator_ac_float_cctor_m_21_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_2_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_3_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_24_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_3_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_72_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_24_nl);
  assign operator_ac_float_cctor_m_21_lpi_1_dfm_1_5_0 = MUX_v_6_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_72_nl,
      6'b111111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_2_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_15_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_14_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_13_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign operator_ac_float_cctor_m_47_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_46_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_47_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_46_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_47_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_69_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_46_nl);
  assign operator_ac_float_cctor_m_47_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_69_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_46_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_21_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_47_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_94_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_21_nl);
  assign operator_ac_float_cctor_m_47_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_94_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_46_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign operator_ac_float_cctor_m_46_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_42_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_43_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_47_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_43_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_70_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_47_nl);
  assign operator_ac_float_cctor_m_46_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_70_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_42_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_22_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_43_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_95_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_22_nl);
  assign operator_ac_float_cctor_m_46_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_95_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_42_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign operator_ac_float_cctor_m_45_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_38_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_39_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_23_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_71_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_not_23_nl);
  assign operator_ac_float_cctor_m_45_lpi_1_dfm_1_5_0 = MUX_v_6_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_71_nl,
      6'b111111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_38_ssc);
  assign operator_ac_float_cctor_m_60_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_38_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_39_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_43_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_43_nl);
  assign operator_ac_float_cctor_m_60_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_38_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_16_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_99_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_not_16_nl);
  assign operator_ac_float_cctor_m_60_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_99_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_38_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_10_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_10_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm);
  assign operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_47_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl = MUX_v_2_2_2(2'b00,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_47_nl);
  assign operator_ac_float_cctor_m_15_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl = MUX_v_4_2_2(4'b0000,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_not_nl);
  assign operator_ac_float_cctor_m_15_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_ssc);
  assign operator_ac_float_cctor_m_30_lpi_1_dfm_1_10_6 = MUX1HOT_v_5_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0,
      5'b01111, 5'b10000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_38_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_39_ssc});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_25_nl = ~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_39_ssc;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_73_nl = MUX_v_6_2_2(6'b000000,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_not_25_nl);
  assign operator_ac_float_cctor_m_30_lpi_1_dfm_1_5_0 = MUX_v_6_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_73_nl,
      6'b111111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_38_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_10_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1_5_0
      = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm);
  assign nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt = conv_s2s_5_6(delay_lane_real_e_0_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[9:5]);
  assign MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt = nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[5:0];
  assign nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt = conv_s2s_5_6(delay_lane_imag_e_1_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[14:10]);
  assign MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt = nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt[5:0];
  assign nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt = conv_s2s_5_6(delay_lane_real_e_1_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[14:10]);
  assign MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt = nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt[5:0];
  assign nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt = conv_s2s_5_6(delay_lane_imag_e_1_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[14:10]);
  assign MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt = nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt[5:0];
  assign nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt = conv_s2s_5_6(delay_lane_real_e_1_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[14:10]);
  assign MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt = nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[5:0];
  assign MAC_9_r_ac_float_2_else_and_nl = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
      & MAC_9_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm;
  assign MAC_9_r_ac_float_2_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2,
      MAC_9_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt
      = conv_s2s_6_7({MAC_9_r_ac_float_2_else_and_nl , MAC_9_r_ac_float_2_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt =
      nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt[6:0];
  assign MAC_10_r_ac_float_3_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4,
      MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign MAC_10_r_ac_float_3_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0,
      MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt
      = conv_s2s_6_7({MAC_10_r_ac_float_3_else_and_nl , MAC_10_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt =
      nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6:0];
  assign MAC_11_r_ac_float_3_else_and_nl = MUX_v_2_2_2(2'b00, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4,
      MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign MAC_11_r_ac_float_3_else_and_1_nl = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0,
      MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt
      = conv_s2s_6_7({MAC_11_r_ac_float_3_else_and_nl , MAC_11_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt =
      nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6:0];
  assign MAC_12_r_ac_float_3_else_and_nl = MUX_v_6_2_2(6'b000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1,
      MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt
      = conv_s2s_6_7(MAC_12_r_ac_float_3_else_and_nl) + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt =
      nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6:0];
  assign MAC_16_r_ac_float_4_else_and_nl = MUX_v_6_2_2(6'b000000, ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1}),
      MAC_16_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt
      = conv_s2s_6_7(MAC_16_r_ac_float_4_else_and_nl) + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt =
      nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6:0];
  assign MAC_9_r_ac_float_3_else_and_nl = operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1
      & MAC_9_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm;
  assign MAC_9_r_ac_float_3_else_and_1_nl = MUX_v_5_2_2(5'b00000, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2,
      MAC_9_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt
      = conv_s2s_6_7({MAC_9_r_ac_float_3_else_and_nl , MAC_9_r_ac_float_3_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt =
      nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6:0];
  assign MAC_9_r_ac_float_4_else_and_nl = operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1
      & MAC_9_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm;
  assign MAC_9_r_ac_float_4_else_and_1_nl = MUX_v_5_2_2(5'b00000, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2,
      MAC_9_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt
      = conv_s2s_6_7({MAC_9_r_ac_float_4_else_and_nl , MAC_9_r_ac_float_4_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt =
      nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_12_cse
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_6_ssc &
      (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_6_cse
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_5_ssc
      & (~ and_dcpl_189);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 = and_1893_cse
      | and_1883_cse;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse = and_1893_cse
      | and_1909_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_1_cse
      = and_2261_cse | and_2264_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_cse
      = ~(and_1909_cse | and_2261_cse | and_2264_cse);
  assign not_tmp_1312 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0!=4'b0000)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4!=2'b00)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6!=5'b00000));
  assign not_tmp_1322 = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0!=4'b0000)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4!=2'b00)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6!=5'b00000));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[4:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_38_nl = ~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_itm
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_38_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[4:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_51_nl = ~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_itm
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_51_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[4:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_53_nl = ~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_itm
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_not_53_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_ssc =
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_8_ssc & (~
      and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_4_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_9_ssc &
      (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_5_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_10_ssc &
      (~ and_dcpl_189);
  assign or_701_nl = and_dcpl_210 | (fsm_output[1]);
  assign mux_433_nl = MUX_s_1_2_2(mux_tmp_146, nor_tmp_6, or_701_nl);
  assign mux_434_nl = MUX_s_1_2_2(mux_433_nl, mux_tmp_380, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_7_ssc = (~(mux_434_nl | (fsm_output[6])))
      | and_dcpl_194;
  assign mux_438_nl = MUX_s_1_2_2(mux_tmp_65, mux_tmp_150, fsm_output[3]);
  assign mux_439_nl = MUX_s_1_2_2(mux_438_nl, mux_tmp_384, fsm_output[2]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_or_8_ssc = (~(mux_439_nl | (fsm_output[6])))
      | and_dcpl_194;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_6_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_2_ssc &
      (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_7_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_3_ssc &
      (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_8_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_5_ssc &
      (~ and_dcpl_189);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_9_ssc
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_7_ssc &
      (~ and_dcpl_189);
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_imag_e_rsci_idat <= 5'b00000;
    end
    else if ( (and_dcpl_169 & ((i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp[5:4]!=2'b01)
        | (~ MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs))
        & and_dcpl_164) | return_imag_e_rsci_idat_mx0c1 ) begin
      return_imag_e_rsci_idat <= MUX_v_5_2_2((i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6[4:0]),
          5'b01111, return_imag_e_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_imag_m_rsci_idat <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_204 ) begin
      return_imag_m_rsci_idat <= MUX1HOT_v_11_3_2(11'b01111111111, 11'b10000000000,
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_itm[12:2]), {i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl
          , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_real_e_rsci_idat <= 5'b00000;
    end
    else if ( (and_dcpl_169 & ((~(MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs
        & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp[4])))
        | (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_l_mux_64_tmp[5]))
        & and_dcpl_164) | return_real_e_rsci_idat_mx0c1 ) begin
      return_real_e_rsci_idat <= MUX_v_5_2_2((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6[4:0]),
          5'b01111, return_real_e_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_real_m_rsci_idat <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_204 ) begin
      return_real_m_rsci_idat <= MUX1HOT_v_11_3_2(11'b01111111111, 11'b10000000000,
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_itm[12:2]), {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl
          , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_or_cse
        ) begin
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl,
          and_dcpl_189);
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_189);
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_189);
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_189);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_nl,
          and_dcpl_189);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_189);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_189);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_189);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_nl,
          and_dcpl_189);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_189);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_189);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_189);
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_nl,
          and_dcpl_189);
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_189);
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_189);
      MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_189);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_197 ) begin
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_16_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_16_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_16_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_15_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_15_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_15_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_15_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_14_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_14_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_14_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_14_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_13_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_13_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_13_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_13_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_6_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5 <= 1'b0;
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4 <= 1'b0;
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0 <= 4'b0000;
      MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_6_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_6_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_5 <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_4 <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0 <= 4'b0000;
      MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5 <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4 <= 1'b0;
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0 <= 4'b0000;
      MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_5_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_3_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_3_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_3_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_3_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_2_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_2_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_2_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_2_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      MAC_1_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= 1'b0;
      MAC_1_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= 1'b0;
      MAC_1_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= 1'b0;
      MAC_1_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= 1'b0;
      reg_return_imag_e_triosy_obj_ld_cse <= 1'b0;
      reg_taps_imag_e_triosy_obj_ld_cse <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= 18'b000000000000000000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0
          <= 4'b0000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0
          <= 4'b0000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0
          <= 4'b0000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0
          <= 4'b0000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_8_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm
          <= 1'b0;
      MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
      MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1
          <= 4'b0000;
    end
    else begin
      MAC_16_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_16_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_16_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_16_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_15_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
      MAC_15_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
      MAC_15_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
      MAC_15_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
      MAC_14_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
      MAC_14_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
      MAC_14_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
      MAC_14_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
      MAC_13_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
      MAC_13_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
      MAC_13_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
      MAC_13_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
      MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_189);
      MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_189);
      MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_189);
      MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_189);
      MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_6_nl,
          and_dcpl_189);
      MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_7_nl,
          and_dcpl_189);
      MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_189);
      MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_189);
      MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_6_nl,
          and_dcpl_189);
      MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_7_nl,
          and_dcpl_189);
      MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_189);
      MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_189);
      MAC_9_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_9_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_9_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_9_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5 <= MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5];
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4 <= MUX1HOT_s_1_19_2((MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[4]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl,
          result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl,
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_1425
          , and_dcpl_1427 , and_dcpl_1428 , and_dcpl_1429 , and_dcpl_1430 , and_dcpl_1431
          , and_dcpl_1432 , and_dcpl_1433 , and_dcpl_1434 , and_dcpl_1435 , and_dcpl_1436
          , and_dcpl_1437 , and_dcpl_1438 , and_dcpl_1439 , and_dcpl_1440});
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0 <= MUX_v_4_2_2(4'b0000,
          mux1h_12_nl, not_1835_nl);
      MAC_6_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_5 <= MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5];
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_4 <= MUX_s_1_2_2((MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[4]),
          (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_conc_32_itm_4_0[4]), and_dcpl_222);
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0 <= MUX1HOT_v_4_10_2((MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[3:0]), (z_out_28[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_108,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_121, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_133,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_138, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_139,
          (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_conc_32_itm_4_0[3:0]),
          {and_dcpl_186 , and_1033_nl , and_1036_nl , and_1039_nl , and_dcpl_192
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_1036 , and_dcpl_222});
      MAC_5_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_5 <= MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5];
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_4 <= MUX_s_1_2_2((MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[4]),
          (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_conc_29_itm_4_0[4]), and_dcpl_222);
      MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0 <= MUX1HOT_v_4_9_2((MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[3:0]),
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1,
          (MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg[3:0]), (z_out[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_107,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_123, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_135,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_137, (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_conc_29_itm_4_0[3:0]),
          {and_dcpl_186 , and_951_nl , and_954_nl , and_957_nl , and_dcpl_192 , and_dcpl_194
          , (~ mux_352_nl) , and_dcpl_198 , and_dcpl_222});
      MAC_5_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
      reg_return_imag_e_triosy_obj_ld_cse <= and_dcpl_223 & and_dcpl_191;
      reg_taps_imag_e_triosy_obj_ld_cse <= ~ or_dcpl_197;
      MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_1_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_1_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_1_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[21:4];
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4
          <= MUX1HOT_v_2_3_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:4]),
          (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0
          <= MUX1HOT_v_4_8_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[3:0]),
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0, (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[3:0]),
          (z_out_1[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_111,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_125, (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          {and_dcpl_186 , and_972_nl , and_975_nl , and_978_nl , and_dcpl_194 , and_dcpl_195
          , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_5_4
          <= MUX1HOT_v_2_3_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:4]),
          (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0
          <= MUX1HOT_v_4_8_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[3:0]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1,
          (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[3:0]), (z_out_29[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_109,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_136, (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          {and_dcpl_186 , and_1043_nl , and_1046_nl , and_1049_nl , and_dcpl_194
          , and_dcpl_195 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_5_4
          <= MUX1HOT_v_2_3_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:4]),
          (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0
          <= MUX1HOT_v_4_8_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[3:0]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2,
          (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[3:0]), (z_out_30[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_124,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_134, (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
          {and_dcpl_186 , and_1150_nl , and_1153_nl , and_1156_nl , and_dcpl_194
          , and_dcpl_195 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_5_4
          <= MUX1HOT_v_2_3_2((MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[5:4]),
          (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0
          <= MUX1HOT_v_4_8_2((MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[3:0]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2,
          (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[3:0]), (z_out_5[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_122,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_132, (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
          {and_dcpl_186 , and_1198_nl , and_1201_nl , and_1204_nl , and_dcpl_194
          , and_dcpl_195 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_5_4
          <= MUX1HOT_v_2_3_2((MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:4]),
          (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5:4]),
          (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0
          <= MUX1HOT_v_4_8_2((MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[3:0]), (z_out_6[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_120,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_130, (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
          (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
          {and_dcpl_186 , and_1243_nl , and_1246_nl , and_1249_nl , and_dcpl_194
          , and_dcpl_195 , and_dcpl_209 , and_dcpl_199});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0
          <= MUX1HOT_v_6_3_2(and_1779_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm[5:0]),
          {(~ mux_184_itm) , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm[6]),
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0
          <= MUX1HOT_v_6_3_2(and_1771_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm[5:0]),
          {(~ mux_184_itm) , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= MUX_v_2_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1[6:5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl,
          and_dcpl_189);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_15_sva_2_1
          <= MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_sva_2_1
          <= MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_15_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva[21]))
          & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_14_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva[21]))
          & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_13_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva[21]))
          & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_12_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva[21]))
          & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_11_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva[21]))
          & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_10_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva[21]))
          & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_8_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva[21]))
          & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_8_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_9_sva[21]))
          & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva[21]))
          & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_7_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_8_sva[21]))
          & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_7_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_8_sva[21]))
          & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva[21]))
          & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_6_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_7_sva[21]))
          & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_6_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_7_sva[21]))
          & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva[21]))
          & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_5_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_6_sva[21]))
          & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_6_sva[21]))
          & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva[21]))
          & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_4_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_5_sva[21]))
          & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva[21]))
          & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_3_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_4_sva[21]))
          & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva[21]))
          & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_2_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_3_sva[21]))
          & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva[21]))
          & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_1_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_2_sva[21]))
          & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva[21]))
          & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
      MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_8_2((~
          MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_102, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_itm_mx0w7,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_194
          , and_dcpl_195 , and_dcpl_198 , and_dcpl_1036});
      MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_8_2((~
          MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          or_897_nl, MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_103, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_1_nl,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_194
          , and_dcpl_195 , and_dcpl_198 , and_dcpl_1036});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_4
          <= MUX1HOT_s_1_18_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_15_nl,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_4,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl,
          result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl,
          {and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_1425 , and_dcpl_1427
          , and_dcpl_1428 , and_dcpl_1429 , and_dcpl_1430 , and_dcpl_1431 , and_dcpl_1432
          , and_dcpl_1433 , and_dcpl_1434 , and_dcpl_1435 , and_dcpl_1436 , and_dcpl_1437
          , and_dcpl_1438 , and_dcpl_1439 , and_dcpl_1440});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0
          <= MUX_v_4_2_2(4'b0000, mux1h_13_nl, not_1837_nl);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_54_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_57_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_60_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_63_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_66_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_69_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_72_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_35_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_38_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_41_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_44_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_47_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_50_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_3[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_53_itm[6]),
          {and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm[5]),
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_107_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm[4:0]),
          operator_ac_float_cctor_e_1_lpi_1_dfm_mx0, operator_ac_float_cctor_e_lpi_1_dfm_mx0,
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm[5]),
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm[5]),
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_0
          <= MUX1HOT_v_5_15_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), operator_ac_float_cctor_m_45_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_60_lpi_1_dfm_1_10_6, (z_out_50[12:8]), (z_out_51[12:8]),
          (z_out_54[12:8]), (z_out_56[12:8]), (z_out_58[12:8]), (z_out_60[12:8]),
          (z_out_61[12:8]), (z_out_64[12:8]), (z_out_65[12:8]), {and_269_itm , and_272_itm
          , and_275_itm , and_278_itm , and_dcpl_277 , and_dcpl_280 , or_dcpl_551
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_1_sva_rsp_1
          <= MUX1HOT_v_6_16_2(MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
          (MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:11]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:11]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:11]), operator_ac_float_cctor_m_45_lpi_1_dfm_1_5_0,
          ({operator_ac_float_cctor_m_60_lpi_1_dfm_1_5_4 , operator_ac_float_cctor_m_60_lpi_1_dfm_1_3_0}),
          (z_out_50[7:2]), (z_out_51[7:2]), (z_out_54[7:2]), (z_out_56[7:2]), (z_out_58[7:2]),
          (z_out_60[7:2]), (z_out_61[7:2]), (z_out_64[7:2]), (z_out_65[7:2]), {and_dcpl_186
          , and_269_itm , and_272_itm , and_275_itm , and_278_itm , and_dcpl_277
          , and_dcpl_280 , or_dcpl_551 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0
          <= MUX1HOT_v_5_22_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_51_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_36_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0, operator_ac_float_cctor_m_63_lpi_1_dfm_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]), (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          operator_ac_float_cctor_m_34_lpi_1_dfm_10_6, operator_i_m_1_lpi_1_dfm_mx0w3_10_6,
          operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0, operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_64_lpi_1_dfm_10_6, operator_ac_float_cctor_m_65_lpi_1_dfm_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
          {and_631_itm , and_634_itm , and_dcpl_596 , and_dcpl_599 , and_636_itm
          , and_640_itm , and_642_itm , nor_270_itm , and_dcpl_195 , and_dcpl_198
          , and_647_itm , nor_286_itm , and_652_itm , and_655_itm , and_660_itm ,
          and_663_itm , and_666_itm , and_670_itm , and_674_itm , and_677_itm , and_680_itm
          , and_684_itm});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_10_6
          <= MUX1HOT_v_5_10_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_36_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_51_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6,
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]), (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          {and_594_ssc , and_597_ssc , and_dcpl_596 , and_dcpl_599 , and_606_ssc
          , and_609_ssc , and_dcpl_552 , and_dcpl_555 , and_dcpl_195 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_5_4
          <= MUX1HOT_v_2_10_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_36_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_51_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4,
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          {and_594_ssc , and_597_ssc , and_dcpl_596 , and_dcpl_599 , and_606_ssc
          , and_609_ssc , and_dcpl_552 , and_dcpl_555 , and_dcpl_195 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_4_sva_3_0
          <= MUX1HOT_v_4_10_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_36_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_51_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0,
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          {and_594_ssc , and_597_ssc , and_dcpl_596 , and_dcpl_599 , and_606_ssc
          , and_609_ssc , and_dcpl_552 , and_dcpl_555 , and_dcpl_195 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0
          <= MUX1HOT_v_2_22_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_51_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_36_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1, operator_ac_float_cctor_m_63_lpi_1_dfm_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0, (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[5:4]),
          operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1, operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_64_lpi_1_dfm_5_4, operator_ac_float_cctor_m_65_lpi_1_dfm_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
          {and_631_itm , and_634_itm , and_dcpl_596 , and_dcpl_599 , and_636_itm
          , and_640_itm , and_642_itm , nor_270_itm , and_dcpl_195 , and_dcpl_198
          , and_647_itm , nor_286_itm , and_652_itm , and_655_itm , and_660_itm ,
          and_663_itm , and_666_itm , and_670_itm , and_674_itm , and_677_itm , and_680_itm
          , and_684_itm});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1
          <= MUX1HOT_v_4_22_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_51_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_36_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2, operator_ac_float_cctor_m_63_lpi_1_dfm_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1, (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[3:0]),
          operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1, operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_64_lpi_1_dfm_3_0, operator_ac_float_cctor_m_65_lpi_1_dfm_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
          {and_631_itm , and_634_itm , and_dcpl_596 , and_dcpl_599 , and_636_itm
          , and_640_itm , and_642_itm , nor_270_itm , and_dcpl_195 , and_dcpl_198
          , and_647_itm , nor_286_itm , and_652_itm , and_655_itm , and_660_itm ,
          and_663_itm , and_666_itm , and_670_itm , and_674_itm , and_677_itm , and_680_itm
          , and_684_itm});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_14_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_14_sva <= delay_lane_imag_e_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_14_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_14_sva <= delay_lane_imag_m_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_14_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_14_sva <= delay_lane_real_e_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_14_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_14_sva <= delay_lane_real_m_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_13_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_13_sva <= delay_lane_imag_e_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_13_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_13_sva <= delay_lane_imag_m_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_13_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_13_sva <= delay_lane_real_e_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_13_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_13_sva <= delay_lane_real_m_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_12_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_12_sva <= delay_lane_imag_e_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_12_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_12_sva <= delay_lane_imag_m_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_12_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_12_sva <= delay_lane_real_e_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_12_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_12_sva <= delay_lane_real_m_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_11_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_11_sva <= delay_lane_imag_e_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_11_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_11_sva <= delay_lane_imag_m_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_11_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_11_sva <= delay_lane_real_e_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_11_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_11_sva <= delay_lane_real_m_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_10_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_10_sva <= delay_lane_imag_e_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_10_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_10_sva <= delay_lane_imag_m_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_10_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_10_sva <= delay_lane_real_e_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_10_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_10_sva <= delay_lane_real_m_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_9_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_9_sva <= delay_lane_imag_e_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_9_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_9_sva <= delay_lane_imag_m_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_9_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_9_sva <= delay_lane_real_e_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_9_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_9_sva <= delay_lane_real_m_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_8_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_8_sva <= delay_lane_imag_e_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_8_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_8_sva <= delay_lane_imag_m_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_8_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_8_sva <= delay_lane_real_e_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_8_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_8_sva <= delay_lane_real_m_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_7_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_7_sva <= delay_lane_imag_e_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_7_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_7_sva <= delay_lane_imag_m_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_7_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_7_sva <= delay_lane_real_e_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_7_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_7_sva <= delay_lane_real_m_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_6_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_6_sva <= delay_lane_imag_e_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_6_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_6_sva <= delay_lane_imag_m_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_6_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_6_sva <= delay_lane_real_e_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_6_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_6_sva <= delay_lane_real_m_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_5_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_5_sva <= delay_lane_imag_e_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_5_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_5_sva <= delay_lane_imag_m_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_5_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_5_sva <= delay_lane_real_e_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_5_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_5_sva <= delay_lane_real_m_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_4_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_4_sva <= delay_lane_imag_e_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_4_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_4_sva <= delay_lane_imag_m_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_4_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_4_sva <= delay_lane_real_e_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_4_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_4_sva <= delay_lane_real_m_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_3_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_3_sva <= delay_lane_imag_e_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_3_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_3_sva <= delay_lane_imag_m_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_3_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_3_sva <= delay_lane_real_e_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_3_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_3_sva <= delay_lane_real_m_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_2_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_2_sva <= delay_lane_imag_e_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_2_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_2_sva <= delay_lane_imag_m_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_2_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_2_sva <= delay_lane_real_e_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_2_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_2_sva <= delay_lane_real_m_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_1_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_1_sva <= delay_lane_imag_e_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_1_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_1_sva <= delay_lane_imag_m_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_1_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_1_sva <= delay_lane_real_e_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_1_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_1_sva <= delay_lane_real_m_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_e_0_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_e_0_sva <= input_imag_e_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_imag_m_0_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_imag_m_0_sva <= input_imag_m_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_e_0_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_e_0_sva <= input_real_e_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_real_m_0_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_197 ) begin
      delay_lane_real_m_0_sva <= input_real_m_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0
          <= 6'b000000;
    end
    else if ( MUX_s_1_2_2(mux_110_nl, mux_109_nl, fsm_output[2]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0
          <= MUX1HOT_v_6_7_2(MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1, z_out_1,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm[5:0]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_199 , and_dcpl_195 , and_dcpl_215
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1
          <= 6'b000000;
    end
    else if ( nor_cse ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0
          <= MUX1HOT_v_6_3_2(and_1827_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm[5:0]),
          {and_dcpl_232 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0
          <= MUX1HOT_v_6_3_2(and_1820_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm[5:0]),
          {and_dcpl_232 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0
          <= MUX1HOT_v_6_3_2(and_1813_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm[5:0]),
          {and_dcpl_232 , and_dcpl_227 , and_dcpl_189});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1
          <= MUX1HOT_v_6_4_2(and_1807_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_63_itm[5:0]),
          {and_dcpl_231 , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1
          <= MUX1HOT_v_6_4_2(and_1801_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_66_itm[5:0]),
          {and_dcpl_231 , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_11_7
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
          <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_11_7
          <= z_out_39[11:7];
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_itm[6]),
          (z_out_39[6]), {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1
          <= MUX1HOT_s_1_4_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_itm[5]),
          (z_out_39[5]), {and_dcpl_186 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1
          <= 6'b000000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7
          <= MUX1HOT_v_5_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6[4:1])), (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[11:7]),
          {and_dcpl_248 , and_dcpl_251 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0
          <= MUX1HOT_s_1_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[6]),
          (operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6[0]), (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[6]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_248 , and_dcpl_251 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1
          <= MUX1HOT_v_6_6_2(and_1791_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_itm[5:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[5:0]),
          ({operator_ac_float_cctor_m_13_lpi_1_dfm_1_5_4 , operator_ac_float_cctor_m_13_lpi_1_dfm_1_3_0}),
          (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[5:0]),
          {and_dcpl_245 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_248 , and_dcpl_251 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_1_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7
          <= MUX1HOT_v_5_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6[4:1])), (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[11:7]),
          {and_dcpl_254 , and_dcpl_257 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0
          <= MUX1HOT_s_1_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[6]),
          (operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6[0]), (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[6]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_254 , and_dcpl_257 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_6_2((and_1787_itm[5:4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_itm[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[5:4]),
          operator_ac_float_cctor_m_7_lpi_1_dfm_1_5_4, (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[5:4]),
          {and_dcpl_245 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_254 , and_dcpl_257 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_6_2((and_1787_itm[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_14_itm[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[3:0]),
          operator_ac_float_cctor_m_7_lpi_1_dfm_1_3_0, (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_sdt[3:0]),
          {and_dcpl_245 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_254 , and_dcpl_257 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_11_7
          <= 5'b00000;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_11_7 <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_1_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_11_7
          <= MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:7];
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_11_7 <= z_out_43[11:7];
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_itm[6]),
          (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[6]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1
          <= MUX1HOT_s_1_4_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_itm[5]),
          (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5]),
          {and_dcpl_186 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2
          <= MUX1HOT_v_5_6_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_3_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_itm[4:0]),
          operator_ac_float_cctor_e_26_lpi_1_dfm_mx0, operator_ac_float_cctor_e_11_lpi_1_dfm_mx0,
          (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[4:0]),
          {and_dcpl_186 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_37_nl
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_38_nl
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_11_7 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_or_2_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_11_7 <= MUX_v_5_2_2((z_out_42[11:7]),
          (z_out_69[11:7]), and_dcpl_215);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_34_lpi_1_dfm_10_6 <= 5'b00000;
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0 <= 2'b00;
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_1_or_ssc ) begin
      operator_ac_float_cctor_m_34_lpi_1_dfm_10_6 <= MUX_v_5_2_2((operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2[10:6]),
          operator_i_m_1_lpi_1_dfm_mx0w3_10_6, and_dcpl_198);
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0 <= MUX1HOT_v_2_3_2((ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0[5:4]),
          (operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2[5:4]), (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[5:4]),
          {and_dcpl_186 , and_dcpl_209 , and_dcpl_198});
      operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1 <= MUX1HOT_v_4_9_2((ac_float_cctor_ac_float_22_2_6_AC_TRN_1_conc_179_itm_5_0[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[3:0]), (z_out_26[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_106,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_119, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_131,
          (operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2[3:0]), (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[3:0]),
          {and_dcpl_186 , and_1135_nl , and_1138_nl , and_1141_nl , and_dcpl_192
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_209 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_2_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_11 <=
          z_out_40[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_3_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_11 <=
          MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_4_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_11 <=
          MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_5_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_11 <=
          MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_6_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_11 <=
          z_out_41[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_11 <=
          1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_7_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_11 <=
          MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_229 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_212 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_6_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_16_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_9_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_15_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[4:0]),
          {and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl
          , and_1469_nl , and_1472_nl , and_1473_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_11_7 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_or_5_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_11_7 <= z_out_44[11:7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_8_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_11_7
          <= MUX1HOT_v_5_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6[4:1])), (z_out_35[11:7]),
          {and_dcpl_367 , and_dcpl_370 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_9_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_11_7
          <= MUX1HOT_v_5_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6[4:1])), (z_out_36[11:7]),
          {and_dcpl_373 , and_dcpl_376 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_10_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_11_7
          <= MUX1HOT_v_5_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6[4:1])), (z_out_37[11:7]),
          {and_dcpl_399 , and_dcpl_402 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_8_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_11_7
          <= MUX1HOT_v_5_3_2((signext_5_4(operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[11:7]),
          (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:7]),
          {and_dcpl_399 , and_dcpl_402 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0
          <= MUX1HOT_s_1_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_itm[6]),
          (operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[6]),
          (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[6]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_399 , and_dcpl_402 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1
          <= MUX1HOT_v_2_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_itm[5:4]),
          operator_ac_float_cctor_m_10_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[5:4]),
          (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_399 , and_dcpl_402 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2
          <= MUX1HOT_v_4_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_itm[3:0]),
          operator_ac_float_cctor_m_10_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[3:0]),
          (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_399 , and_dcpl_402 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_ssc )
        begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), operator_ac_float_cctor_m_39_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_54_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_5_4 <=
          MUX1HOT_v_2_4_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), operator_ac_float_cctor_m_39_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_54_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_3_0 <=
          MUX1HOT_v_4_4_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), operator_ac_float_cctor_m_39_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_54_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6
          <= MUX1HOT_v_5_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_57_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_42_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_65_lpi_1_dfm_10_6,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0, operator_r_m_8_lpi_1_dfm_mx0w6_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4
          <= MUX1HOT_v_2_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_57_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_42_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_65_lpi_1_dfm_5_4,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1, operator_r_m_8_lpi_1_dfm_mx0w6_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0
          <= MUX1HOT_v_4_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_57_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_42_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_65_lpi_1_dfm_3_0,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1, operator_r_m_8_lpi_1_dfm_mx0w6_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_1_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6
          <= MUX1HOT_v_5_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_43_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_58_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_65_lpi_1_dfm_10_6, operator_r_m_9_lpi_1_dfm_mx0w6_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4
          <= MUX1HOT_v_2_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_43_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_58_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_65_lpi_1_dfm_5_4, operator_r_m_9_lpi_1_dfm_mx0w6_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0
          <= MUX1HOT_v_4_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_43_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_58_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_65_lpi_1_dfm_3_0, operator_r_m_9_lpi_1_dfm_mx0w6_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_484 , and_dcpl_487 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_4_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6
          <= MUX1HOT_v_5_5_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2[10:6]),
          operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_10_6, operator_r_m_1_lpi_1_dfm_mx0w4_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4 <=
          MUX1HOT_v_2_5_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2[5:4]),
          operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_5_4, (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[5:4]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0 <=
          MUX1HOT_v_4_5_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_29_lpi_1_dfm_mx0w2[3:0]),
          operator_ac_float_cctor_m_19_lpi_1_dfm_mx0w3_3_0, (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[3:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_3_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_37_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_52_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_5_4
          <= MUX1HOT_v_2_4_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_37_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_52_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_3_0
          <= MUX1HOT_v_4_4_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_37_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_52_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_5_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_4_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_52_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_37_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_5_4
          <= MUX1HOT_v_2_4_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_52_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_37_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_3_0
          <= MUX1HOT_v_4_4_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_52_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_37_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_6_sva_mx0c1
          , and_dcpl_689 , and_dcpl_692});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_5_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_38_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_53_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_5_4
          <= MUX1HOT_v_2_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_38_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_53_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_3_0
          <= MUX1HOT_v_4_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_38_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_53_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_7_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_6_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_53_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_38_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_5_4
          <= MUX1HOT_v_2_4_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_53_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_38_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_3_0
          <= MUX1HOT_v_4_4_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_53_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_38_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_8_sva_mx0c1
          , and_dcpl_854 , and_dcpl_857});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= 1'b0;
    end
    else if ( (~(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg)) | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva[21])
        | (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= ~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4 <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_ssc )
        begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4 <= ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_1_nl
          & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_8_ssc);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0 <=
          MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_28_nl,
          4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_8_ssc);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_9_sva[21]) | (~
        MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg & (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_9_sva
          <= ~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c4
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg,
          MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[4:0]),
          5'b01111, {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva[21]) | (~(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= ~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c4
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c5
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c6
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c7
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva <= MUX1HOT_v_5_8_2(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_4_lpi_1_dfm_1_4_0,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_4_lpi_1_dfm_1_5_0[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0,
          operator_ac_float_cctor_e_19_lpi_1_dfm, operator_ac_float_cctor_e_65_lpi_1_dfm,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[4:0]),
          {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_9_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_5_nl ,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_7_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c4
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c5
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c6});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva[21]) | (~(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_10_sva
          <= ~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c4
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg,
          MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[4:0]),
          5'b01111, {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva[21]) | (~(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= ~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4 <=
          1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_2_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_4 <=
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_5_nl &
          (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_10_ssc);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_3_0 <=
          MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_18_nl,
          4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_10_ssc);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva[21]) |
        (~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg & (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_11_sva
          <= ~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva[21]) | (~(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= ~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c4
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c5
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c6
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c7
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c8
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva <= MUX1HOT_v_5_9_2(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_5_lpi_1_dfm_1_4_0,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_5_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_10_lpi_1_dfm_1_5_0[4:0]),
          operator_ac_float_cctor_e_3_lpi_1_dfm, operator_ac_float_cctor_e_29_lpi_1_dfm,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[4:0]),
          {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_11_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_17_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_19_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_21_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_23_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c5
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c6
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c7});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva[21]) |
        (~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg & (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_12_sva
          <= ~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva[21]) | (~(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= ~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4 <=
          1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_1_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4 <=
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_3_nl &
          (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c6);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0 <=
          ~(MUX_v_4_2_2(nor_566_nl, 4'b1111, or_1068_nl));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c4
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c5
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c6
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c7
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c8
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva <= MUX1HOT_v_5_9_2(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_6_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_6_lpi_1_dfm_1_5_0[4:0]),
          operator_ac_float_cctor_e_31_lpi_1_dfm, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1_5_0[4:0]),
          operator_ac_float_cctor_e_33_lpi_1_dfm, operator_ac_float_cctor_e_14_lpi_1_dfm,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[4:0]),
          {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_12_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_25_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_27_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_29_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c5
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c6
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c7});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva[21]) |
        (~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg & (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_13_sva
          <= ~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= 1'b0;
    end
    else if ( (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
        | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva[21]) | (~(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
        & MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= ~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4 <=
          1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_5_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4 <=
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_11_nl
          & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_13_ssc);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0 <=
          MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_29_nl,
          4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_13_ssc);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_14_sva[21]) |
        (~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg & (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_14_sva
          <= ~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_8_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), operator_ac_float_cctor_m_54_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_39_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_5_4
          <= MUX1HOT_v_2_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), operator_ac_float_cctor_m_54_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_39_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_3_0
          <= MUX1HOT_v_4_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), operator_ac_float_cctor_m_54_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_39_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_sva_mx0c1
          , and_dcpl_452 , and_dcpl_455});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_15_sva_2_1
          <= MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c4
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c5
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c6
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva <= MUX1HOT_v_5_7_2(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_8_lpi_1_dfm_1_5_0[4:0]),
          operator_ac_float_cctor_e_29_lpi_1_dfm, operator_ac_float_cctor_e_14_lpi_1_dfm,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[4:0]),
          {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_14_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_37_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_39_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c4
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c5});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_15_sva[21]) |
        (~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg & (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_15_sva
          <= ~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1
          <= 2'b00;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_sva_2_1
          <= MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva <= 5'b00000;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c4
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg,
          MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[4:0]),
          5'b01111, {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva
          <= 1'b0;
    end
    else if ( (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_sva[21]) | (~
        MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm)
        | (~(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg & (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])))
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_sva
          <= ~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_15_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_sva[21]))
          & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_15_sva[21]))
          & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_13_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_14_sva[21]))
          & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva[21]))
          & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_12_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva[21]))
          & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva[21]))
          & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva[21]))
          & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva[21]))
          & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm
          <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_195 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_nl,
          my_complex_float_t_cctor_imag_operator_return_4_sva_mx0w1, and_dcpl_195);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva[21]))
          & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nand_9_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva[21]))
          & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva[21]))
          & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm
          <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_212 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_nl,
          my_complex_float_t_cctor_real_operator_return_9_sva_mx0w1, and_dcpl_212);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_257 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= ~(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva[21]))
          & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_29_sva <= 1'b0;
      ac_float_cctor_operator_return_12_sva <= 1'b0;
      ac_float_cctor_operator_return_17_sva <= 1'b0;
      ac_float_cctor_operator_return_42_sva <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_cse
        ) begin
      ac_float_cctor_operator_return_29_sva <= MUX1HOT_s_1_4_2((~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_11_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl, ac_float_cctor_operator_return_2_sva_mx0w2,
          MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      ac_float_cctor_operator_return_12_sva <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_7_nl,
          ac_float_cctor_operator_return_12_sva_mx0w1, ac_float_cctor_operator_return_16_sva_mx0w2,
          my_complex_float_t_cctor_imag_operator_return_14_sva_mx0w2, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      ac_float_cctor_operator_return_17_sva <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_8_nl,
          ac_float_cctor_operator_return_27_sva_mx0w1, ac_float_cctor_operator_return_17_sva_mx0w2,
          my_complex_float_t_cctor_imag_operator_return_sva_mx0w6, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      ac_float_cctor_operator_return_42_sva <= MUX1HOT_s_1_4_2((~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          ac_float_cctor_operator_return_42_sva_mx0w1, ac_float_cctor_operator_return_47_sva_mx0w2,
          my_complex_float_t_cctor_real_operator_return_9_sva_mx0w1, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_3_sva <= 1'b0;
      ac_float_cctor_operator_return_31_sva <= 1'b0;
      ac_float_cctor_operator_return_32_sva <= 1'b0;
      ac_float_cctor_operator_return_59_sva <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_cse
        ) begin
      ac_float_cctor_operator_return_3_sva <= MUX1HOT_s_1_3_2((~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_16_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_operator_return_31_sva <= MUX1HOT_s_1_3_2((~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_13_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl, my_complex_float_t_cctor_imag_operator_return_4_sva_mx0w1,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_operator_return_32_sva <= MUX1HOT_s_1_3_2((~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_14_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl, my_complex_float_t_cctor_imag_operator_return_13_sva_mx0w2,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_operator_return_59_sva <= MUX1HOT_s_1_3_2((~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_11_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, my_complex_float_t_cctor_imag_operator_return_14_sva_mx0w2,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_30_sva <= 1'b0;
      ac_float_cctor_operator_return_48_sva <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_zero_or_1_cse
        ) begin
      ac_float_cctor_operator_return_30_sva <= MUX1HOT_s_1_4_2((~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_12_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl, ac_float_cctor_operator_return_46_sva_mx0w2,
          my_complex_float_t_cctor_imag_operator_return_3_sva_mx0w3, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_operator_return_48_sva <= MUX1HOT_s_1_4_2((~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1),
          ac_float_cctor_operator_return_57_sva_mx0w1, ac_float_cctor_operator_return_48_sva_mx0w2,
          MAC_10_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_60_sva <= 1'b0;
      ac_float_cctor_operator_return_61_sva <= 1'b0;
      ac_float_cctor_operator_return_62_sva <= 1'b0;
      ac_float_cctor_operator_return_63_sva <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_op2_zero_or_2_cse
        ) begin
      ac_float_cctor_operator_return_60_sva <= MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_1_nl,
          MAC_12_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, MAC_11_my_complex_float_t_cctor_imag_operator_my_complex_float_t_cctor_imag_operator_nor_tmp,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_198});
      ac_float_cctor_operator_return_61_sva <= MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_2_nl,
          MAC_13_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, my_complex_float_t_cctor_imag_operator_return_3_sva_mx0w3,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_198});
      ac_float_cctor_operator_return_62_sva <= MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_3_nl,
          MAC_14_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, my_complex_float_t_cctor_imag_operator_return_4_sva_mx0w1,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_198});
      ac_float_cctor_operator_return_63_sva <= MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_4_nl,
          MAC_15_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl, my_complex_float_t_cctor_imag_operator_return_13_sva_mx0w2,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_dcpl_192 | and_dcpl_194
        | and_dcpl_195 | and_dcpl_212 ) begin
      MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_7_2((~
          MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl,
          my_complex_float_t_cctor_imag_operator_return_sva_mx0w6, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_194 , and_dcpl_195
          , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_dcpl_192 | and_dcpl_194
        | and_dcpl_195 | and_dcpl_198 ) begin
      MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_7_2((~
          MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          or_899_nl, MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl,
          my_complex_float_t_cctor_real_operator_return_10_sva_mx0w6, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , and_dcpl_194 , and_dcpl_195
          , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
      MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_1_cse )
        begin
      MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_6_2((~
          MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl,
          my_complex_float_t_cctor_real_operator_return_10_sva_mx0w6, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_212});
      MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_6_2((~
          MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl,
          my_complex_float_t_cctor_real_operator_return_11_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_212});
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_6_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_1_nl,
          MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_itm_mx0w7,
          my_complex_float_t_cctor_real_operator_return_12_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_212});
      MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_6_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_10_nl,
          MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl,
          my_complex_float_t_cctor_real_operator_return_4_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_199 | and_dcpl_194 | and_dcpl_195
        ) begin
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_5_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_11_nl,
          MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl,
          my_complex_float_t_cctor_imag_operator_return_3_sva_mx0w3, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
      MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
      MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_3_cse ) begin
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_6_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_12_nl,
          MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl,
          my_complex_float_t_cctor_real_operator_return_11_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_198});
      MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_6_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_13_nl,
          MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl,
          my_complex_float_t_cctor_real_operator_return_12_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_198});
      MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_6_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_2_nl,
          MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl,
          my_complex_float_t_cctor_real_operator_return_4_sva_mx0w5, {and_dcpl_189
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_194 , and_dcpl_195 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
    end
    else if ( and_dcpl_189 | and_dcpl_209 | and_dcpl_194 | and_dcpl_195 | and_dcpl_198
        ) begin
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_5_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_3_nl,
          or_898_nl, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_9_nl,
          MAC_6_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_194 , and_dcpl_195 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= 1'b0;
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= 1'b0;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_4_cse ) begin
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_4_nl,
          MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl,
          MAC_7_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_194 , and_dcpl_198});
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_5_nl,
          MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl,
          MAC_8_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_194 , and_dcpl_198});
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_6_nl,
          MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl,
          MAC_9_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl,
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_194 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_14_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c3 | operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c4
        ) begin
      operator_ac_float_cctor_e_14_lpi_1_dfm <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c3 , operator_ac_float_cctor_e_14_lpi_1_dfm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_19_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c3 | operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c4
        ) begin
      operator_ac_float_cctor_e_19_lpi_1_dfm <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_9_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c3 , operator_ac_float_cctor_e_19_lpi_1_dfm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_29_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c3 | operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c4
        ) begin
      operator_ac_float_cctor_e_29_lpi_1_dfm <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_9_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c3 , operator_ac_float_cctor_e_29_lpi_1_dfm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_3_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_3_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_3_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_31_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c3 | operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c4
        ) begin
      operator_ac_float_cctor_e_31_lpi_1_dfm <= MUX1HOT_v_5_5_2(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_11_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_13_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c3 , operator_ac_float_cctor_e_31_lpi_1_dfm_mx0c4});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_33_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_33_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_13_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_33_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_34_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_34_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_14_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_34_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_61_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_61_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_11_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_61_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_62_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_62_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_12_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_62_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_63_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_63_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_13_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_63_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_64_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_64_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_14_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_64_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_e_65_lpi_1_dfm <= 5'b00000;
    end
    else if ( and_dcpl_189 | operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c1 | operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c2
        | operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c3 ) begin
      operator_ac_float_cctor_e_65_lpi_1_dfm <= MUX1HOT_v_5_4_2(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_15_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[4:0]),
          {and_dcpl_189 , operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c1 , operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c2
          , operator_ac_float_cctor_e_65_lpi_1_dfm_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0 <= 5'b00000;
    end
    else if ( ((~(mux_443_nl | (fsm_output[6]))) | and_dcpl_192) & (and_dcpl_189
        | and_dcpl_209 | and_dcpl_199 | and_969_rgt | or_487_rgt) ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0 <= MUX1HOT_v_5_6_2(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg,
          MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[4:0]),
          5'b01111, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_mx0w1[4:0]),
          {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_969_rgt , operator_13_2_true_AC_TRN_AC_WRAP_1_and_16_nl
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_11_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4 <= operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_6_nl
          & (~ operator_13_2_true_AC_TRN_AC_WRAP_1_and_21_ssc);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0 <= MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_13_nl,
          4'b1111, operator_13_2_true_AC_TRN_AC_WRAP_1_and_21_ssc);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6 <= 5'b00000;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_7_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6 <= MUX1HOT_v_5_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          operator_r_m_4_lpi_1_dfm_mx0w5_10_6, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1[10:6]),
          {and_462_ssc , and_465_ssc , and_468_ssc , and_471_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4 <= MUX1HOT_v_2_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          operator_r_m_4_lpi_1_dfm_mx0w5_5_4, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1[5:4]),
          {and_462_ssc , and_465_ssc , and_468_ssc , and_471_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0 <= MUX1HOT_v_4_7_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          operator_r_m_4_lpi_1_dfm_mx0w5_3_0, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_mx0w1[3:0]),
          {and_462_ssc , and_465_ssc , and_468_ssc , and_471_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6 <= 5'b00000;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_8_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6 <= MUX1HOT_v_5_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          operator_r_m_14_lpi_1_dfm_mx0w5_10_6, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[10:6]),
          {and_506_ssc , and_509_ssc , and_512_ssc , and_515_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4 <= MUX1HOT_v_2_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          operator_r_m_14_lpi_1_dfm_mx0w5_5_4, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[5:4]),
          {and_506_ssc , and_509_ssc , and_512_ssc , and_515_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0 <= MUX1HOT_v_4_7_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          operator_r_m_14_lpi_1_dfm_mx0w5_3_0, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[3:0]),
          {and_506_ssc , and_509_ssc , and_512_ssc , and_515_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6 <= 5'b00000;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_10_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6 <= MUX1HOT_v_5_6_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), operator_r_m_7_lpi_1_dfm_mx0w4_10_6,
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[10:6]), {and_581_ssc
          , and_584_ssc , and_587_ssc , and_590_ssc , and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4 <= MUX1HOT_v_2_6_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), operator_r_m_7_lpi_1_dfm_mx0w4_5_4,
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[5:4]), {and_581_ssc
          , and_584_ssc , and_587_ssc , and_590_ssc , and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0 <= MUX1HOT_v_4_6_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), operator_r_m_7_lpi_1_dfm_mx0w4_3_0,
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[3:0]), {and_581_ssc
          , and_584_ssc , and_587_ssc , and_590_ssc , and_dcpl_198 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
          <= 6'b000000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_6_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_11_6
          <= MUX1HOT_v_6_7_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[11:6]),
          ({{1{operator_ac_float_cctor_m_lpi_1_dfm_1_10_6[4]}}, operator_ac_float_cctor_m_lpi_1_dfm_1_10_6}),
          ({{1{operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6[4]}}, operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6}),
          (z_out_35[11:6]), (z_out_33[11:6]), ({{1{ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6[4]}},
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6}),
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[11:6]),
          {and_dcpl_361 , and_dcpl_364 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_420
          , and_dcpl_423 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_5_4
          <= MUX1HOT_v_2_7_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[5:4]),
          operator_ac_float_cctor_m_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_17_lpi_1_dfm_1_5_4,
          (z_out_35[5:4]), (z_out_33[5:4]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4,
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {and_dcpl_361 , and_dcpl_364 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_420
          , and_dcpl_423 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_26_itm_3_0
          <= MUX1HOT_v_4_7_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[3:0]),
          operator_ac_float_cctor_m_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_17_lpi_1_dfm_1_3_0,
          (z_out_35[3:0]), (z_out_33[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0,
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {and_dcpl_361 , and_dcpl_364 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_420
          , and_dcpl_423 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6
          <= 6'b000000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_7_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6
          <= MUX1HOT_v_6_5_2(({{1{operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6[4]}},
          operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6}), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[11:6]),
          (z_out_35[11:6]), ({{1{operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6[4]}},
          operator_ac_float_cctor_m_17_lpi_1_dfm_1_10_6}), (z_out_39[11:6]), {and_dcpl_432
          , and_dcpl_435 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4
          <= MUX1HOT_v_2_5_2(operator_ac_float_cctor_m_20_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[5:4]),
          (z_out_35[5:4]), operator_ac_float_cctor_m_17_lpi_1_dfm_1_5_4, (z_out_39[5:4]),
          {and_dcpl_432 , and_dcpl_435 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0
          <= MUX1HOT_v_4_5_2(operator_ac_float_cctor_m_20_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[3:0]),
          (z_out_35[3:0]), operator_ac_float_cctor_m_17_lpi_1_dfm_1_3_0, (z_out_39[3:0]),
          {and_dcpl_432 , and_dcpl_435 , and_dcpl_1575 , and_dcpl_1578 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva <= z_out_45;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva <= z_out_46;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva <= z_out_47;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva <= z_out_42;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva <= z_out_43;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva <= z_out_44;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
          <= nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva[1:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= 2'b00;
    end
    else if ( and_dcpl_199 | and_dcpl_195 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= MUX_v_2_2_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0,
          MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl,
          and_dcpl_195);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva <= MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_rshift_itm;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_486 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
          <= r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0 <= 1'b0;
    end
    else if ( ~ or_dcpl_486 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0 <= z_out_48[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0 <=
          1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0 <=
          1'b0;
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva
          <= 2'b00;
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= 2'b00;
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva
          <= 2'b00;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_8_cse
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0 <=
          MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_16_sva_1[0]),
          (z_out_49[0]), and_dcpl_194);
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0 <=
          MUX_s_1_2_2((z_out_49[0]), (z_out_48[0]), and_dcpl_194);
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva
          <= MUX_v_2_2_2(MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0,
          and_dcpl_194);
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= MUX_v_2_2_2(MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0,
          and_dcpl_194);
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva
          <= MUX_v_2_2_2(MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0,
          and_dcpl_194);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 2'b00;
    end
    else if ( and_dcpl_199 | and_dcpl_194 | and_dcpl_215 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= MUX1HOT_v_2_3_2(MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0,
          {and_dcpl_199 , and_dcpl_194 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_507 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva <= z_out_46;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_507 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva <= z_out_45;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva <= 13'b0000000000000;
    end
    else if ( ~ or_dcpl_507 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva <= z_out_47;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva
          <= r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0 <=
          1'b0;
    end
    else if ( ~ or_dcpl_507 ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0 <=
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_mx0w0[0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_507 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva
          <= 2'b00;
    end
    else if ( and_dcpl_192 | and_dcpl_195 | and_dcpl_215 ) begin
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva
          <= MUX1HOT_v_2_3_2(i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_mx0w0,
          MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva_mx0w0,
          {and_dcpl_192 , and_dcpl_195 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_509 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva
          <= 2'b00;
    end
    else if ( ~ or_dcpl_509 ) begin
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva
          <= i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_or_ssc )
        begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0
          <= ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_1_nl
          & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c6)
          & (~ or_dcpl_558);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1
          <= ~(MUX_v_4_2_2(nor_574_nl, 4'b1111, or_dcpl_558));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1
          <= 6'b000000;
    end
    else if ( ~((~ mux_128_nl) | and_dcpl_189) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1, (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_194 , and_dcpl_215 , and_dcpl_227});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_0
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1
          <= 6'b000000;
    end
    else if ( reg_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_1_cse
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1
          <= MUX1HOT_v_6_4_2(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          z_out_28, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1,
          (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_194 , and_dcpl_227});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1
          <= MUX1HOT_v_6_4_2(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
          z_out_30, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1,
          (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_194 , and_dcpl_227});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1
          <= MUX1HOT_v_6_4_2(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
          z_out_29, i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1,
          (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_194 , and_dcpl_227});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_0
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_0
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1
          <= 6'b000000;
    end
    else if ( ~((mux_130_nl & and_dcpl_206) | and_dcpl_189) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1
          <= MUX1HOT_v_6_4_2(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1, z_out, (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_195 , and_dcpl_227});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_0
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1
          <= 6'b000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_or_5_cse )
        begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_54_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_2_sva_mx0w1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_57_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_60_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          z_out_2, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_44_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_47_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
          z_out_3, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_50_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_95_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~(mux_551_nl | (fsm_output[6:4]!=3'b000)) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1
          <= MUX1HOT_v_6_4_2(and_1795_nl, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_69_itm[5:0]),
          {and_236_nl , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1
          <= MUX1HOT_v_6_6_2(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          z_out_2, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_20_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_72_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_195 , and_dcpl_227 , and_dcpl_189
          , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1
          <= MUX1HOT_v_6_6_2(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_21_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_35_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_195 , and_dcpl_227 , and_dcpl_189
          , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1
          <= MUX1HOT_v_6_6_2(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_22_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_38_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_195 , and_dcpl_227 , and_dcpl_189
          , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1
          <= MUX1HOT_v_6_6_2(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
          r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_23_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_41_itm[5:0]),
          {and_dcpl_186 , and_dcpl_199 , and_dcpl_195 , and_dcpl_227 , and_dcpl_189
          , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_195 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1
          <= MUX1HOT_v_6_5_2(MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
          i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_3[5:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_53_itm[5:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_90_cse , and_dcpl_194
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_195 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[5]),
          (z_out_3[5]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm[5]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_90_cse , and_dcpl_194
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_195 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1
          <= MUX1HOT_v_5_6_2((MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[4:0]),
          (z_out_3[4:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm[4:0]),
          MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_and_90_cse , and_dcpl_194
          , and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_71_cse
          , and_dcpl_199});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt[5]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[5]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm[5]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_sdt[4:0]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[4:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm[4:0]),
          MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt[5]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[5]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm[5]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_sdt[4:0]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[4:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm[4:0]),
          MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt[5]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm[5]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_203 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_sdt[4:0]),
          (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[4:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm[4:0]),
          MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_82_cse , and_dcpl_199
          , and_dcpl_227 , and_dcpl_189 , and_dcpl_209});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_194 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[5]),
          (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm[5]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( ~ and_dcpl_194 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1
          <= MUX1HOT_v_5_6_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_sdt[4:0]),
          (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[4:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm[4:0]),
          MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl,
          MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_cse , and_dcpl_192
          , and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_71_cse
          , and_dcpl_199});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc
        & (or_736_rgt | and_1462_rgt | and_1465_rgt | and_1466_rgt) ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2
          <= MUX1HOT_v_5_8_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_conc_57_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_and_15_itm[4:0]),
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_qr_6_0_12_lpi_1_dfm_1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_14_lpi_1_dfm_1_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[4:0]),
          (z_out_39[4:0]), {and_dcpl_186 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_33_nl
          , and_1462_rgt , and_1465_rgt , and_1466_rgt , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_33_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_0 <= MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt[6]),
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3[6]), and_dcpl_194);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_1 <= MUX1HOT_s_1_3_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0[5]),
          (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt[5]),
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3[5]), {and_dcpl_186
          , and_dcpl_243 , and_dcpl_194});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_0 <= MUX1HOT_s_1_4_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0[4]),
          (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt[4]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_8_nl, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3[4]),
          {and_dcpl_186 , and_dcpl_243 , (~ mux_119_itm) , and_dcpl_194});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1 <= MUX1HOT_v_4_4_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_31_itm_5_0[3:0]),
          (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_sdt[3:0]),
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_1_nl, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_mx0w3[3:0]),
          {and_dcpl_186 , and_dcpl_243 , (~ mux_119_itm) , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( (mux_553_nl | (~(nor_536_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_6))
        | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_itm
        & (fsm_output[1:0]==2'b11)))) & nor_774_cse & and_dcpl_184 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_109_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_itm[4:0]),
          operator_ac_float_cctor_e_23_lpi_1_dfm_mx0, operator_ac_float_cctor_e_8_lpi_1_dfm_mx0,
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1
          <= 5'b00000;
    end
    else if ( (mux_555_nl | (~(nor_534_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_6))
        | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
        & (fsm_output[1:0]==2'b11)))) & nor_774_cse & and_dcpl_184 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm_5_0_rsp_1
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_111_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_itm[4:0]),
          operator_ac_float_cctor_e_24_lpi_1_dfm_mx0, operator_ac_float_cctor_e_9_lpi_1_dfm_mx0,
          {and_dcpl_186 , and_dcpl_227 , and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_35_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0 <= MUX1HOT_s_1_4_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6]),
          (z_out_68[6]), (z_out_69[6]), (z_out_70[6]), {and_dcpl_243 , and_dcpl_199
          , and_dcpl_194 , and_dcpl_215});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1 <= MUX1HOT_s_1_5_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0[5]),
          (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[5]),
          (z_out_68[5]), (z_out_69[5]), (z_out_70[5]), {and_dcpl_186 , and_dcpl_243
          , and_dcpl_199 , and_dcpl_194 , and_dcpl_215});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2 <= MUX1HOT_v_5_7_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_34_itm_5_0[4:0]),
          (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[4:0]),
          operator_ac_float_cctor_e_27_lpi_1_dfm_mx0, operator_ac_float_cctor_e_12_lpi_1_dfm_mx0,
          (z_out_68[4:0]), (z_out_69[4:0]), (z_out_70[4:0]), {and_dcpl_186 , and_dcpl_243
          , operator_13_2_true_AC_TRN_AC_WRAP_1_and_22_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_23_nl
          , and_dcpl_199 , and_dcpl_194 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_38_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0 <= MUX1HOT_s_1_3_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6]),
          (z_out_42[6]), (z_out_69[6]), {and_dcpl_243 , and_dcpl_192 , and_dcpl_215});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1 <= MUX1HOT_s_1_4_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0[5]),
          (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[5]),
          (z_out_42[5]), (z_out_69[5]), {and_dcpl_186 , and_dcpl_243 , and_dcpl_192
          , and_dcpl_215});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2 <= MUX1HOT_v_5_6_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_37_itm_5_0[4:0]),
          (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[4:0]),
          operator_ac_float_cctor_e_28_lpi_1_dfm_mx0, operator_ac_float_cctor_e_13_lpi_1_dfm_mx0,
          (z_out_42[4:0]), (z_out_69[4:0]), {and_dcpl_186 , and_dcpl_243 , operator_13_2_true_AC_TRN_AC_WRAP_1_and_24_nl
          , operator_13_2_true_AC_TRN_AC_WRAP_1_and_25_nl , and_dcpl_192 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_41_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0 <= MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6]),
          (z_out_43[6]), and_dcpl_192);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1 <= MUX1HOT_s_1_3_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0[5]),
          (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[5]),
          (z_out_43[5]), {and_dcpl_186 , and_dcpl_243 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2 <= MUX1HOT_v_5_5_2((operator_13_2_true_AC_TRN_AC_WRAP_1_conc_40_itm_5_0[4:0]),
          (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[4:0]),
          operator_ac_float_cctor_e_21_lpi_1_dfm_mx0, ({operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_4
          , operator_ac_float_cctor_e_6_lpi_1_dfm_mx0_3_0}), (z_out_43[4:0]), {and_dcpl_186
          , and_dcpl_243 , operator_13_2_true_AC_TRN_AC_WRAP_1_and_26_nl , operator_13_2_true_AC_TRN_AC_WRAP_1_and_27_nl
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1
          <= MUX_v_6_2_2(and_1765_nl, (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[5:0]),
          and_dcpl_227);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1
          <= 6'b000000;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1
          <= MUX_v_6_2_2(and_1759_nl, (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[5:0]),
          and_dcpl_227);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0 <= 5'b00000;
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1 <= 2'b00;
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_ssc ) begin
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0 <= MUX1HOT_v_5_3_2((operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2[10:6]),
          operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_10_6, operator_r_m_1_lpi_1_dfm_mx0w4_10_6,
          {and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1 <= MUX1HOT_v_2_4_2((ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0[5:4]),
          (operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2[5:4]), operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_5_4,
          (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[5:4]), {and_dcpl_186 , and_dcpl_209
          , and_dcpl_199 , and_dcpl_198});
      operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2 <= MUX1HOT_v_4_10_2((ac_float_cctor_ac_float_22_2_6_AC_TRN_2_conc_176_itm_5_0[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[3:0]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_105, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_117,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_129, (operator_ac_float_cctor_m_44_lpi_1_dfm_mx0w2[3:0]),
          operator_ac_float_cctor_m_49_lpi_1_dfm_mx0w3_3_0, (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[3:0]),
          {and_dcpl_186 , and_1184_nl , and_1187_nl , and_1190_nl , and_dcpl_192
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0
          <= 5'b00000;
    end
    else if ( MUX_s_1_2_2(mux_557_nl, nor_789_nl, or_6_cse) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0
          <= MUX1HOT_v_5_15_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_60_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_45_lpi_1_dfm_1_10_6, (z_out_53[12:8]), (z_out_52[12:8]),
          (z_out_66[12:8]), (z_out_67[12:8]), (z_out_63[12:8]), (z_out_59[12:8]),
          (z_out_57[12:8]), (z_out_62[12:8]), (z_out_55[12:8]), {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c4
          , and_dcpl_277 , and_dcpl_280 , or_dcpl_551 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1
          <= 6'b000000;
    end
    else if ( and_dcpl_186 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c3
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c4
        | and_dcpl_277 | and_dcpl_280 | and_dcpl_194 | and_dcpl_195 | and_dcpl_198
        | and_dcpl_212 | and_dcpl_282 | and_dcpl_285 | and_dcpl_286 | and_dcpl_287
        | and_dcpl_288 | and_dcpl_291 | and_dcpl_292 | and_dcpl_293 | and_dcpl_294
        | and_dcpl_296 | and_dcpl_297 | and_dcpl_298 | and_dcpl_299 | and_dcpl_300
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1
          <= MUX1HOT_v_6_16_2(MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
          (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:11]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:11]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:11]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:11]), ({operator_ac_float_cctor_m_60_lpi_1_dfm_1_5_4
          , operator_ac_float_cctor_m_60_lpi_1_dfm_1_3_0}), operator_ac_float_cctor_m_45_lpi_1_dfm_1_5_0,
          (z_out_53[7:2]), (z_out_52[7:2]), (z_out_66[7:2]), (z_out_67[7:2]), (z_out_63[7:2]),
          (z_out_59[7:2]), (z_out_57[7:2]), (z_out_62[7:2]), (z_out_55[7:2]), {and_dcpl_186
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_mx0c4
          , and_dcpl_277 , and_dcpl_280 , or_dcpl_551 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_10_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_14_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_18_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_22_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_26_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_30_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_34_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_38_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0
          <= 5'b00000;
    end
    else if ( mux_562_nl & nor_796_cse ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0
          <= MUX1HOT_v_5_10_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_46_lpi_1_dfm_1_10_6, (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]), (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          operator_i_m_8_lpi_1_dfm_mx0w10_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4
          , and_dcpl_327 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0
          <= 5'b00000;
    end
    else if ( mux_566_nl & nor_796_cse ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0
          <= MUX1HOT_v_5_10_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_47_lpi_1_dfm_1_10_6, (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]), (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          operator_i_m_9_lpi_1_dfm_mx0w10_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4
          , and_dcpl_345 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_26_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0
          <= MUX1HOT_v_5_8_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]), operator_r_m_2_lpi_1_dfm_mx0w6_10_6,
          (z_out_40[10:6]), {and_568_itm , and_571_itm , and_574_itm , and_577_itm
          , and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_9_2((MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:4]),
          (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]), operator_r_m_2_lpi_1_dfm_mx0w6_5_4,
          (z_out_40[5:4]), {and_dcpl_186 , and_568_itm , and_571_itm , and_574_itm
          , and_577_itm , and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_9_2((MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[3:0]),
          (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]), operator_r_m_2_lpi_1_dfm_mx0w6_3_0,
          (z_out_40[3:0]), {and_dcpl_186 , and_568_itm , and_571_itm , and_574_itm
          , and_577_itm , and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_27_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0
          <= MUX1HOT_v_5_8_2((MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]), operator_r_m_3_lpi_1_dfm_mx0w6_10_6,
          (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[10:6]),
          {and_618_itm , and_621_itm , and_624_itm , and_627_itm , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_9_2((MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:4]),
          (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]), operator_r_m_3_lpi_1_dfm_mx0w6_5_4,
          (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {and_dcpl_186 , and_618_itm , and_621_itm , and_624_itm , and_627_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_9_2((MAC_7_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[3:0]),
          (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]), operator_r_m_3_lpi_1_dfm_mx0w6_3_0,
          (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {and_dcpl_186 , and_618_itm , and_621_itm , and_624_itm , and_627_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_28_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0
          <= MUX1HOT_v_5_8_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]), operator_r_m_4_lpi_1_dfm_mx0w5_10_6,
          (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[10:6]),
          {and_705_itm , and_708_itm , and_711_itm , and_714_itm , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_9_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[5:4]),
          (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]), operator_r_m_4_lpi_1_dfm_mx0w5_5_4,
          (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {and_dcpl_186 , and_705_itm , and_708_itm , and_711_itm , and_714_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_9_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_itm[3:0]),
          (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]), operator_r_m_4_lpi_1_dfm_mx0w5_3_0,
          (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {and_dcpl_186 , and_705_itm , and_708_itm , and_711_itm , and_714_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_29_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0
          <= MUX1HOT_v_5_8_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[12:8]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]), operator_r_m_14_lpi_1_dfm_mx0w5_10_6,
          (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[10:6]),
          {and_784_itm , and_787_itm , and_790_itm , and_793_itm , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_9_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[5:4]),
          (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), operator_r_m_14_lpi_1_dfm_mx0w5_5_4,
          (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {and_dcpl_186 , and_784_itm , and_787_itm , and_790_itm , and_793_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_9_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[3:0]),
          (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), operator_r_m_14_lpi_1_dfm_mx0w5_3_0,
          (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {and_dcpl_186 , and_784_itm , and_787_itm , and_790_itm , and_793_itm ,
          and_dcpl_195 , and_dcpl_198 , and_dcpl_212 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_30_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0
          <= MUX1HOT_v_5_6_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_r_m_15_lpi_1_dfm_mx0w4_10_6,
          (z_out_41[10:6]), {and_870_itm , and_873_itm , and_876_itm , and_879_itm
          , and_dcpl_195 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_7_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[5:4]),
          (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_r_m_15_lpi_1_dfm_mx0w4_5_4,
          (z_out_41[5:4]), {and_dcpl_186 , and_870_itm , and_873_itm , and_876_itm
          , and_879_itm , and_dcpl_195 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_7_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm[3:0]),
          (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_r_m_15_lpi_1_dfm_mx0w4_3_0,
          (z_out_41[3:0]), {and_dcpl_186 , and_870_itm , and_873_itm , and_876_itm
          , and_879_itm , and_dcpl_195 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_31_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0
          <= MUX1HOT_v_5_7_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[21:17]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[21:17]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          operator_r_m_3_lpi_1_dfm_mx0w6_10_6, (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[10:6]),
          {and_1318_itm , and_1321_itm , and_1324_itm , and_1327_itm , and_dcpl_195
          , and_dcpl_198 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0
          <= MUX1HOT_v_2_8_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[5:4]),
          (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          operator_r_m_3_lpi_1_dfm_mx0w6_5_4, (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[5:4]),
          {and_dcpl_186 , and_1318_itm , and_1321_itm , and_1324_itm , and_1327_itm
          , and_dcpl_195 , and_dcpl_198 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1
          <= MUX1HOT_v_4_8_2((MAC_8_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_itm[3:0]),
          (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          operator_r_m_3_lpi_1_dfm_mx0w6_3_0, (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_sdt[3:0]),
          {and_dcpl_186 , and_1318_itm , and_1321_itm , and_1324_itm , and_1327_itm
          , and_dcpl_195 , and_dcpl_198 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1 <= 6'b000000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_44_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_0 <= MUX_s_1_2_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6]),
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_mx0w2[6]), and_dcpl_192);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1 <= MUX1HOT_v_6_5_2(MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
          MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp,
          MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp,
          (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[5:0]),
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_mx0w2[5:0]), {and_dcpl_186
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_243 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0 <=
          2'b00;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_0 <=
          MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6:5];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1 <=
          5'b00000;
    end
    else if ( ~ and_dcpl_189 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1 <=
          MUX1HOT_v_5_3_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[4:0]),
          operator_ac_float_cctor_e_25_lpi_1_dfm_mx0, operator_ac_float_cctor_e_10_lpi_1_dfm_mx0,
          {and_dcpl_227 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1 <= 5'b00000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_46_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0 <= MUX_v_2_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[6:5]),
          (z_out_44[6:5]), and_dcpl_192);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1 <= MUX1HOT_v_5_6_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_sdt[4:0]),
          operator_ac_float_cctor_e_22_lpi_1_dfm_mx0, operator_ac_float_cctor_e_7_lpi_1_dfm_mx0,
          operator_ac_float_cctor_e_30_lpi_1_dfm_mx0, operator_ac_float_cctor_e_15_lpi_1_dfm_mx0,
          (z_out_44[4:0]), {and_dcpl_243 , and_1537_nl , and_1541_nl , and_1544_nl
          , and_1548_nl , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_48_cse ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_0 <= MUX_v_2_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6:5]),
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2[6:5]), and_dcpl_192);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4 <= MUX1HOT_s_1_4_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[4]),
          operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_4, operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_4,
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2[4]), {and_dcpl_243
          , operator_13_2_true_AC_TRN_AC_WRAP_1_and_31_ssc , operator_13_2_true_AC_TRN_AC_WRAP_1_and_32_ssc
          , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0 <= MUX1HOT_v_4_4_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[3:0]),
          operator_ac_float_cctor_e_35_lpi_1_dfm_mx0_3_0, operator_ac_float_cctor_e_20_lpi_1_dfm_mx0_3_0,
          (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2[3:0]), {and_dcpl_243
          , operator_13_2_true_AC_TRN_AC_WRAP_1_and_31_ssc , operator_13_2_true_AC_TRN_AC_WRAP_1_and_32_ssc
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_2_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_0
          <= MUX1HOT_v_5_5_2((signext_5_4(operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[11:7]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          (z_out_38[11:7]), (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          {and_dcpl_254 , and_dcpl_257 , and_dcpl_199 , and_dcpl_194 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_3_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_0
          <= MUX1HOT_v_5_5_2((signext_5_4(operator_ac_float_cctor_m_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[11:7]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          (z_out_35[11:7]), (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          {and_dcpl_361 , and_dcpl_364 , and_dcpl_199 , and_dcpl_194 , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_4_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_0
          <= MUX1HOT_v_5_4_2((signext_5_4(operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[11:7]),
          (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          (z_out_33[11:7]), {and_dcpl_367 , and_dcpl_370 , and_dcpl_199 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_6_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_itm[6]),
          (operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[6]),
          (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          (z_out_33[6]), {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_367 , and_dcpl_370 , and_dcpl_199 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1
          <= MUX1HOT_v_2_6_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_itm[5:4]),
          operator_ac_float_cctor_m_8_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[5:4]),
          (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:4]),
          (z_out_33[5:4]), {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_367 , and_dcpl_370 , and_dcpl_199 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2
          <= MUX1HOT_v_4_6_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_and_itm[3:0]),
          operator_ac_float_cctor_m_8_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[3:0]),
          (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          (z_out_33[3:0]), {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse
          , and_dcpl_189 , and_dcpl_367 , and_dcpl_370 , and_dcpl_199 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_5_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_0
          <= MUX1HOT_v_5_4_2((signext_5_4(operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[11:7]),
          (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          {and_dcpl_373 , and_dcpl_376 , and_dcpl_199 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_6_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_0
          <= MUX1HOT_v_5_6_2((signext_5_4(operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6[4:1])), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[11:7]),
          (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          (MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          {and_dcpl_379 , and_dcpl_382 , and_dcpl_385 , and_dcpl_388 , and_dcpl_192
          , and_dcpl_195});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_or_7_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_0
          <= MUX1HOT_v_5_4_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6[4:1])), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          (MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:7]),
          {and_dcpl_392 , and_dcpl_395 , and_dcpl_192 , and_dcpl_195});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
          <= 5'b00000;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_0
          <= MUX1HOT_v_5_6_2((signext_5_4(operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[11:7]),
          (signext_5_4(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[4:1])),
          (z_out_33[11:7]), (z_out_34[11:7]), (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          {and_dcpl_405 , and_dcpl_408 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_6
          <= MUX1HOT_s_1_8_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl,
          (operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[0]),
          (z_out_33[6]), (z_out_34[6]), (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_405 , and_dcpl_408 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_0
          <= MUX1HOT_v_2_8_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_itm[5:4]),
          operator_ac_float_cctor_m_6_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[5:4]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4,
          (z_out_33[5:4]), (z_out_34[5:4]), (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_405 , and_dcpl_408 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_rsp_1_5_0_rsp_1
          <= MUX1HOT_v_4_8_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_itm[3:0]),
          operator_ac_float_cctor_m_6_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[3:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0,
          (z_out_33[3:0]), (z_out_34[3:0]), (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_cse ,
          and_dcpl_189 , and_dcpl_405 , and_dcpl_408 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_1_itm_mx0c5
          , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6[4:1])), (signext_5_4(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6[4:1])),
          (z_out_33[11:7]), (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          {and_dcpl_379 , and_dcpl_382 , and_dcpl_420 , and_dcpl_423 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6
          <= MUX1HOT_s_1_6_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[6]),
          (operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6[0]),
          (z_out_33[6]), (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_420 , and_dcpl_423
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4
          <= MUX1HOT_v_2_6_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[5:4]),
          operator_ac_float_cctor_m_11_lpi_1_dfm_1_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4,
          (z_out_33[5:4]), (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_420 , and_dcpl_423
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0
          <= MUX1HOT_v_4_6_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[3:0]),
          operator_ac_float_cctor_m_11_lpi_1_dfm_1_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0,
          (z_out_33[3:0]), (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_420 , and_dcpl_423
          , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_2_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0
          <= MUX1HOT_v_5_5_2((signext_5_4(operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[11:7]),
          (z_out_34[11:7]), (signext_5_4(operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6[4:1])),
          (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[11:7]),
          {and_dcpl_392 , and_dcpl_395 , and_dcpl_426 , and_dcpl_429 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6
          <= MUX1HOT_s_1_6_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6]),
          (operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[6]),
          (z_out_34[6]), (operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6[0]), (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4
          <= MUX1HOT_v_2_6_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[5:4]),
          operator_ac_float_cctor_m_12_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[5:4]),
          (z_out_34[5:4]), operator_ac_float_cctor_m_16_lpi_1_dfm_1_5_4, (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0
          <= MUX1HOT_v_4_6_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[3:0]),
          operator_ac_float_cctor_m_12_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[3:0]),
          (z_out_34[3:0]), operator_ac_float_cctor_m_16_lpi_1_dfm_1_3_0, (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_3_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_0
          <= MUX1HOT_v_5_5_2((signext_5_4(operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6[4:1])),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6[4:1])), (z_out_34[11:7]),
          (z_out_38[11:7]), {and_dcpl_248 , and_dcpl_251 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_2_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6
          <= MUX1HOT_s_1_6_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6]),
          (operator_ac_float_cctor_m_13_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[6]),
          (operator_ac_float_cctor_m_16_lpi_1_dfm_1_10_6[0]), (z_out_34[6]), (z_out_38[6]),
          {and_dcpl_243 , and_dcpl_248 , and_dcpl_251 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0
          <= MUX1HOT_v_2_6_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[5:4]),
          operator_ac_float_cctor_m_13_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[5:4]),
          operator_ac_float_cctor_m_16_lpi_1_dfm_1_5_4, (z_out_34[5:4]), (z_out_38[5:4]),
          {and_dcpl_243 , and_dcpl_248 , and_dcpl_251 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1
          <= MUX1HOT_v_4_6_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[3:0]),
          operator_ac_float_cctor_m_13_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_9_sva_1[3:0]),
          operator_ac_float_cctor_m_16_lpi_1_dfm_1_3_0, (z_out_34[3:0]), (z_out_38[3:0]),
          {and_dcpl_243 , and_dcpl_248 , and_dcpl_251 , and_dcpl_426 , and_dcpl_429
          , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_4_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_0
          <= MUX1HOT_v_5_6_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6[4:1])), (z_out_33[11:7]),
          (signext_5_4(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[4:1])),
          (z_out_34[11:7]), (z_out_41[11:7]), {and_dcpl_432 , and_dcpl_435 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
          , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_3_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6
          <= MUX1HOT_s_1_7_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[6]),
          (operator_ac_float_cctor_m_20_lpi_1_dfm_1_10_6[0]), (z_out_33[6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6[0]),
          (z_out_34[6]), (z_out_41[6]), {and_dcpl_243 , and_dcpl_432 , and_dcpl_435
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0
          <= MUX1HOT_v_2_7_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[5:4]),
          operator_ac_float_cctor_m_20_lpi_1_dfm_1_5_4, (z_out_33[5:4]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4,
          (z_out_34[5:4]), (z_out_41[5:4]), {and_dcpl_243 , and_dcpl_432 , and_dcpl_435
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
          , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1
          <= MUX1HOT_v_4_7_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_16_sva_1[3:0]),
          operator_ac_float_cctor_m_20_lpi_1_dfm_1_3_0, (z_out_33[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0,
          (z_out_34[3:0]), (z_out_41[3:0]), {and_dcpl_243 , and_dcpl_432 , and_dcpl_435
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c3
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c4
          , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_mx0c5
          , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0
          <= 5'b00000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_5_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6[4:1])), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[11:7]),
          (signext_5_4(operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6[4:1])), (z_out_40[11:7]),
          {and_dcpl_405 , and_dcpl_408 , and_dcpl_385 , and_dcpl_388 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0
          <= 5'b00000;
    end
    else if ( MUX_s_1_2_2(mux_569_nl, nor_809_nl, or_6_cse) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_0
          <= MUX1HOT_v_5_22_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_41_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_56_lpi_1_dfm_1_10_6, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6,
          operator_ac_float_cctor_m_63_lpi_1_dfm_10_6, (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]), operator_i_m_1_lpi_1_dfm_mx0w3_10_6,
          operator_ac_float_cctor_m_34_lpi_1_dfm_10_6, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0, operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0,
          operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0, operator_ac_float_cctor_m_64_lpi_1_dfm_10_6,
          operator_ac_float_cctor_m_65_lpi_1_dfm_10_6, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5
          , and_dcpl_195 , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1 <= 4'b0000;
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0 <= 5'b00000;
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1 <= 2'b00;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_2_or_1_ssc ) begin
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1 <= MUX1HOT_v_4_8_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2,
          (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[3:0]), (z_out_19[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_118,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_128, (operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1[3:0]),
          operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_3_0, operator_r_m_15_lpi_1_dfm_mx0w4_3_0,
          {and_1285_nl , and_1288_nl , and_1291_nl , and_dcpl_194 , and_dcpl_195
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_0 <= MUX1HOT_v_5_3_2((operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1[10:6]),
          operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_10_6, operator_r_m_15_lpi_1_dfm_mx0w4_10_6,
          {and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
      operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1 <= MUX1HOT_v_2_3_2((operator_ac_float_cctor_m_59_lpi_1_dfm_mx0w1[5:4]),
          operator_ac_float_cctor_m_50_lpi_1_dfm_mx0w2_5_4, operator_r_m_15_lpi_1_dfm_mx0w4_5_4,
          {and_dcpl_209 , and_dcpl_199 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1 <= 4'b0000;
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0 <= 5'b00000;
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1 <= 2'b00;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_6_ssc ) begin
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1 <= MUX1HOT_v_4_7_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[3:0]), (z_out_22[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_116,
          (operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1[3:0]), operator_ac_float_cctor_m_46_lpi_1_dfm_1_3_0,
          operator_r_m_lpi_1_dfm_mx0w6_3_0, {and_1334_nl , and_1337_nl , and_1340_nl
          , and_dcpl_194 , and_dcpl_209 , and_dcpl_327 , and_dcpl_198});
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_0 <= MUX1HOT_v_5_3_2((operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1[10:6]),
          operator_ac_float_cctor_m_46_lpi_1_dfm_1_10_6, operator_r_m_lpi_1_dfm_mx0w6_10_6,
          {and_dcpl_209 , and_dcpl_327 , and_dcpl_198});
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1 <= MUX1HOT_v_2_3_2((operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1[5:4]),
          operator_ac_float_cctor_m_46_lpi_1_dfm_1_5_4, operator_r_m_lpi_1_dfm_mx0w6_5_4,
          {and_dcpl_209 , and_dcpl_327 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1 <= 4'b0000;
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0 <= 5'b00000;
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1 <= 2'b00;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_7_ssc ) begin
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1 <= MUX1HOT_v_4_7_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg[3:0]), (z_out_3[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_114,
          (operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1[3:0]), operator_ac_float_cctor_m_47_lpi_1_dfm_1_3_0,
          operator_i_m_6_lpi_1_dfm_mx0w4_3_0, {and_942_nl , and_945_nl , and_948_nl
          , and_dcpl_194 , and_dcpl_209 , and_dcpl_345 , and_dcpl_198});
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_0 <= MUX1HOT_v_5_3_2((operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1[10:6]),
          operator_ac_float_cctor_m_47_lpi_1_dfm_1_10_6, operator_i_m_6_lpi_1_dfm_mx0w4_10_6,
          {and_dcpl_209 , and_dcpl_345 , and_dcpl_198});
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1 <= MUX1HOT_v_2_3_2((operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1[5:4]),
          operator_ac_float_cctor_m_47_lpi_1_dfm_1_5_4, operator_i_m_6_lpi_1_dfm_mx0w4_5_4,
          {and_dcpl_209 , and_dcpl_345 , and_dcpl_198});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_1_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), operator_ac_float_cctor_m_40_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_55_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_5_4 <=
          MUX1HOT_v_2_4_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), operator_ac_float_cctor_m_40_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_55_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_3_0 <=
          MUX1HOT_v_4_4_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), operator_ac_float_cctor_m_40_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_55_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_2_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_2_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), operator_ac_float_cctor_m_55_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_40_lpi_1_dfm_1_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4 <=
          MUX1HOT_v_2_4_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), operator_ac_float_cctor_m_55_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_40_lpi_1_dfm_1_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0 <=
          MUX1HOT_v_4_4_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), operator_ac_float_cctor_m_55_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_40_lpi_1_dfm_1_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_mx0c1
          , and_dcpl_496 , and_dcpl_499});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_or_2_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6
          <= MUX1HOT_v_5_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[21:17]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[21:17]), operator_ac_float_cctor_m_58_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_43_lpi_1_dfm_1_10_6, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6,
          operator_r_m_lpi_1_dfm_mx0w6_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_552 , and_dcpl_555 , and_dcpl_195});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4
          <= MUX1HOT_v_2_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[16:15]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[16:15]), operator_ac_float_cctor_m_58_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_43_lpi_1_dfm_1_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4,
          operator_r_m_lpi_1_dfm_mx0w6_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_552 , and_dcpl_555 , and_dcpl_195});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0
          <= MUX1HOT_v_4_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_rshift_itm[14:11]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_3_lshift_itm[14:11]), operator_ac_float_cctor_m_58_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_43_lpi_1_dfm_1_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0,
          operator_r_m_lpi_1_dfm_mx0w6_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_mx0c1
          , and_dcpl_521 , and_dcpl_524 , and_dcpl_552 , and_dcpl_555 , and_dcpl_195});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_3_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_10_6
          <= MUX1HOT_v_5_5_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2[10:6]),
          operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_10_6, operator_i_m_1_lpi_1_dfm_mx0w3_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4 <=
          MUX1HOT_v_2_5_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2[5:4]),
          operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_5_4, (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[5:4]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0 <=
          MUX1HOT_v_4_5_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_14_lpi_1_dfm_mx0w2[3:0]),
          operator_ac_float_cctor_m_18_lpi_1_dfm_mx0w3_3_0, (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[3:0]),
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_5_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6
          <= MUX1HOT_v_5_5_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2[10:6]),
          operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_10_6, operator_r_m_15_lpi_1_dfm_mx0w4_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4 <=
          MUX1HOT_v_2_5_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2[5:4]),
          operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_5_4, operator_r_m_15_lpi_1_dfm_mx0w4_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0 <=
          MUX1HOT_v_4_5_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2[3:0]),
          operator_ac_float_cctor_m_2_lpi_1_dfm_mx0w3_3_0, operator_r_m_15_lpi_1_dfm_mx0w4_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_6_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_10_6
          <= MUX1HOT_v_5_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2[10:6]),
          operator_r_m_lpi_1_dfm_mx0w6_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4 <=
          MUX1HOT_v_2_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2[5:4]),
          operator_r_m_lpi_1_dfm_mx0w6_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0 <=
          MUX1HOT_v_4_4_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2[3:0]),
          operator_r_m_lpi_1_dfm_mx0w6_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_1_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6
          <= MUX1HOT_v_5_22_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_56_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_41_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_64_lpi_1_dfm_10_6,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0, operator_r_m_2_lpi_1_dfm_mx0w6_10_6,
          operator_r_m_1_lpi_1_dfm_mx0w4_10_6, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , and_dcpl_799 , and_dcpl_802 , and_dcpl_198
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4
          <= MUX1HOT_v_2_22_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_56_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_41_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_64_lpi_1_dfm_5_4,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1, operator_r_m_2_lpi_1_dfm_mx0w6_5_4,
          (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[5:4]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , and_dcpl_799 , and_dcpl_802 , and_dcpl_198
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0
          <= MUX1HOT_v_4_22_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_56_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_41_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_64_lpi_1_dfm_3_0,
          operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2, operator_r_m_2_lpi_1_dfm_mx0w6_3_0,
          (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[3:0]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , and_dcpl_799 , and_dcpl_802 , and_dcpl_198
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c7
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_mx0c21});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_7_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6
          <= MUX1HOT_v_5_5_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2[10:6]),
          operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_10_6, operator_i_m_6_lpi_1_dfm_mx0w4_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4 <=
          MUX1HOT_v_2_5_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2[5:4]),
          operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_5_4, operator_i_m_6_lpi_1_dfm_mx0w4_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0 <=
          MUX1HOT_v_4_5_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2[3:0]),
          operator_ac_float_cctor_m_48_lpi_1_dfm_mx0w3_3_0, operator_i_m_6_lpi_1_dfm_mx0w4_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_mx0c1
          , and_dcpl_209 , and_dcpl_199 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6
          <= 5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_2_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_10_6
          <= MUX1HOT_v_5_24_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), operator_ac_float_cctor_m_42_lpi_1_dfm_1_10_6,
          operator_ac_float_cctor_m_57_lpi_1_dfm_1_10_6, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_0,
          operator_ac_float_cctor_m_64_lpi_1_dfm_10_6, (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]), operator_r_m_1_lpi_1_dfm_mx0w4_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_10_6,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_10_6, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_10_6,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_10_6,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_799 , and_dcpl_802 , and_dcpl_195
          , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_5_4
          <= MUX1HOT_v_2_24_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_42_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_57_lpi_1_dfm_1_5_4, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_64_lpi_1_dfm_5_4, (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[5:4]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_5_4,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_5_4, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_5_4,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_799 , and_dcpl_802 , and_dcpl_195
          , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_3_0
          <= MUX1HOT_v_4_24_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_42_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_57_lpi_1_dfm_1_3_0, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2,
          operator_ac_float_cctor_m_64_lpi_1_dfm_3_0, (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (operator_r_m_1_lpi_1_dfm_mx0w4_5_0[3:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_7_sva_3_0,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_7_sva_10_0_rsp_1_rsp_1,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0,
          operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_2_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_3_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_4_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_5_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_6_sva_10_0_rsp_1_rsp_1,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c1
          , and_dcpl_478 , and_dcpl_481 , and_dcpl_799 , and_dcpl_802 , and_dcpl_195
          , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c21
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c22
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_8_sva_mx0c23});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6 <=
          5'b00000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4 <=
          2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0 <=
          4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_or_9_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6 <=
          MUX1HOT_v_5_4_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2[10:6]),
          operator_i_m_7_lpi_1_dfm_mx0w3_10_6, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4 <=
          MUX1HOT_v_2_4_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2[5:4]),
          operator_i_m_7_lpi_1_dfm_mx0w3_5_4, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0 <=
          MUX1HOT_v_4_4_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2[3:0]),
          operator_i_m_7_lpi_1_dfm_mx0w3_3_0, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
          , and_dcpl_209 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6 <= 5'b00000;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_and_9_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_10_6 <= MUX1HOT_v_5_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[21:17]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[21:17]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:17]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:17]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:8]),
          operator_r_m_6_lpi_1_dfm_mx0w5_10_6, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1[10:6]),
          {and_537_ssc , and_540_ssc , and_543_ssc , and_546_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_5_4 <= MUX1HOT_v_2_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[16:15]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[16:15]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          operator_r_m_6_lpi_1_dfm_mx0w5_5_4, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1[5:4]),
          {and_537_ssc , and_540_ssc , and_543_ssc , and_546_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0 <= MUX1HOT_v_4_7_2((MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[14:11]),
          (MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[14:11]), (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          operator_r_m_6_lpi_1_dfm_mx0w5_3_0, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_mx0w1[3:0]),
          {and_537_ssc , and_540_ssc , and_543_ssc , and_546_ssc , and_dcpl_195 ,
          and_dcpl_198 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_ac_float_cctor_m_65_lpi_1_dfm_10_6 <= 5'b00000;
      operator_ac_float_cctor_m_65_lpi_1_dfm_5_4 <= 2'b00;
      operator_ac_float_cctor_m_65_lpi_1_dfm_3_0 <= 4'b0000;
      operator_ac_float_cctor_m_64_lpi_1_dfm_10_6 <= 5'b00000;
      operator_ac_float_cctor_m_64_lpi_1_dfm_5_4 <= 2'b00;
      operator_ac_float_cctor_m_64_lpi_1_dfm_3_0 <= 4'b0000;
      operator_ac_float_cctor_m_63_lpi_1_dfm_10_6 <= 5'b00000;
      operator_ac_float_cctor_m_63_lpi_1_dfm_5_4 <= 2'b00;
      operator_ac_float_cctor_m_63_lpi_1_dfm_3_0 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_3_or_8_cse ) begin
      operator_ac_float_cctor_m_65_lpi_1_dfm_10_6 <= MUX_v_5_2_2((operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0[10:6]),
          operator_i_m_9_lpi_1_dfm_mx0w10_10_6, and_dcpl_198);
      operator_ac_float_cctor_m_65_lpi_1_dfm_5_4 <= MUX_v_2_2_2((operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0[5:4]),
          operator_i_m_9_lpi_1_dfm_mx0w10_5_4, and_dcpl_198);
      operator_ac_float_cctor_m_65_lpi_1_dfm_3_0 <= MUX_v_4_2_2((operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0[3:0]),
          operator_i_m_9_lpi_1_dfm_mx0w10_3_0, and_dcpl_198);
      operator_ac_float_cctor_m_64_lpi_1_dfm_10_6 <= MUX_v_5_2_2((operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0[10:6]),
          operator_i_m_8_lpi_1_dfm_mx0w10_10_6, and_dcpl_198);
      operator_ac_float_cctor_m_64_lpi_1_dfm_5_4 <= MUX_v_2_2_2((operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0[5:4]),
          operator_i_m_8_lpi_1_dfm_mx0w10_5_4, and_dcpl_198);
      operator_ac_float_cctor_m_64_lpi_1_dfm_3_0 <= MUX_v_4_2_2((operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0[3:0]),
          operator_i_m_8_lpi_1_dfm_mx0w10_3_0, and_dcpl_198);
      operator_ac_float_cctor_m_63_lpi_1_dfm_10_6 <= MUX_v_5_2_2((operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0[10:6]),
          operator_i_m_7_lpi_1_dfm_mx0w3_10_6, and_dcpl_198);
      operator_ac_float_cctor_m_63_lpi_1_dfm_5_4 <= MUX_v_2_2_2((operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0[5:4]),
          operator_i_m_7_lpi_1_dfm_mx0w3_5_4, and_dcpl_198);
      operator_ac_float_cctor_m_63_lpi_1_dfm_3_0 <= MUX_v_4_2_2((operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0[3:0]),
          operator_i_m_7_lpi_1_dfm_mx0w3_3_0, and_dcpl_198);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_1_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0
          <= MUX1HOT_v_2_11_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0[5:4]),
          (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_46_lpi_1_dfm_1_5_4, (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]), (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          operator_i_m_8_lpi_1_dfm_mx0w10_5_4, {and_dcpl_186 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4
          , and_dcpl_327 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1
          <= MUX1HOT_v_4_11_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_23_itm_5_0[3:0]),
          (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_46_lpi_1_dfm_1_3_0, (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]), (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          operator_i_m_8_lpi_1_dfm_mx0w10_3_0, {and_dcpl_186 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c4
          , and_dcpl_327 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_or_2_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0
          <= MUX1HOT_v_2_11_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0[5:4]),
          (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[16:15]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[16:15]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_47_lpi_1_dfm_1_5_4, (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]), (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[7:6]),
          operator_i_m_9_lpi_1_dfm_mx0w10_5_4, {and_dcpl_186 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4
          , and_dcpl_345 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1
          <= MUX1HOT_v_4_11_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_conc_24_itm_5_0[3:0]),
          (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_rshift_itm[14:11]),
          (MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_1_lshift_itm[14:11]), (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_47_lpi_1_dfm_1_3_0, (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]), (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_1_lshift_itm[5:2]),
          operator_i_m_9_lpi_1_dfm_mx0w10_3_0, {and_dcpl_186 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c3
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c4
          , and_dcpl_345 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_mx0c6
          , and_dcpl_194 , and_dcpl_195 , and_dcpl_198 , and_dcpl_212});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_12_cse
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_7_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[6]),
          (operator_ac_float_cctor_m_11_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[6]),
          (operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[6]),
          (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          (MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_385 , and_dcpl_388
          , and_dcpl_192 , and_dcpl_195});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_0
          <= MUX1HOT_v_2_7_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[5:4]),
          operator_ac_float_cctor_m_11_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[5:4]),
          operator_ac_float_cctor_m_15_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[5:4]),
          (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          (MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:4]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_385 , and_dcpl_388
          , and_dcpl_192 , and_dcpl_195});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1
          <= MUX1HOT_v_4_7_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_sdt[3:0]),
          operator_ac_float_cctor_m_11_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_7_sva_1[3:0]),
          operator_ac_float_cctor_m_15_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[3:0]),
          (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          (MAC_1_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          {and_dcpl_243 , and_dcpl_379 , and_dcpl_382 , and_dcpl_385 , and_dcpl_388
          , and_dcpl_192 , and_dcpl_195});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_6_cse
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0
          <= MUX1HOT_s_1_6_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[6]),
          (operator_ac_float_cctor_m_6_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[6]),
          (operator_ac_float_cctor_m_15_lpi_1_dfm_1_10_6[0]), (z_out_40[6]), {and_dcpl_243
          , and_dcpl_405 , and_dcpl_408 , and_dcpl_385 , and_dcpl_388 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0
          <= MUX1HOT_v_2_6_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[5:4]),
          operator_ac_float_cctor_m_6_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[5:4]),
          operator_ac_float_cctor_m_15_lpi_1_dfm_1_5_4, (z_out_40[5:4]), {and_dcpl_243
          , and_dcpl_405 , and_dcpl_408 , and_dcpl_385 , and_dcpl_388 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1
          <= MUX1HOT_v_4_6_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_sdt[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_2_sva_1[3:0]),
          operator_ac_float_cctor_m_6_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_11_sva_1[3:0]),
          operator_ac_float_cctor_m_15_lpi_1_dfm_1_3_0, (z_out_40[3:0]), {and_dcpl_243
          , and_dcpl_405 , and_dcpl_408 , and_dcpl_385 , and_dcpl_388 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1
          <= 4'b0000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_or_ssc
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_0
          <= MUX1HOT_v_2_22_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[16:15]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[16:15]), operator_ac_float_cctor_m_41_lpi_1_dfm_1_5_4,
          operator_ac_float_cctor_m_56_lpi_1_dfm_1_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4,
          operator_ac_float_cctor_m_63_lpi_1_dfm_5_4, (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[5:4]),
          operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_0_rsp_1, operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_0_rsp_1,
          operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_0_rsp_1, operator_ac_float_cctor_m_64_lpi_1_dfm_5_4,
          operator_ac_float_cctor_m_65_lpi_1_dfm_5_4, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5
          , and_dcpl_195 , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_rsp_1_rsp_1
          <= MUX1HOT_v_4_22_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_rshift_itm[14:11]),
          (MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_2_lshift_itm[14:11]), operator_ac_float_cctor_m_41_lpi_1_dfm_1_3_0,
          operator_ac_float_cctor_m_56_lpi_1_dfm_1_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0,
          operator_ac_float_cctor_m_63_lpi_1_dfm_3_0, (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (operator_i_m_1_lpi_1_dfm_mx0w3_5_0[3:0]),
          operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1, operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2,
          operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1, operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1,
          operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1, operator_ac_float_cctor_m_64_lpi_1_dfm_3_0,
          operator_ac_float_cctor_m_65_lpi_1_dfm_3_0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c1
          , and_dcpl_720 , and_dcpl_723 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c4
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c5
          , and_dcpl_195 , and_dcpl_198 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c8
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c9
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c10
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c11
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c12
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c13
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c14
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c15
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c16
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c17
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c18
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c19
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c20
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_6_sva_mx0c21});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[6]),
          (operator_ac_float_cctor_m_8_lpi_1_dfm_1_10_6[0]), (z_out_35[6]), {and_dcpl_243
          , and_dcpl_367 , and_dcpl_370 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_1
          <= MUX1HOT_v_2_4_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[5:4]),
          operator_ac_float_cctor_m_8_lpi_1_dfm_1_5_4, (z_out_35[5:4]), {and_dcpl_243
          , and_dcpl_367 , and_dcpl_370 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2
          <= MUX1HOT_v_4_4_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_4_sva_1[3:0]),
          operator_ac_float_cctor_m_8_lpi_1_dfm_1_3_0, (z_out_35[3:0]), {and_dcpl_243
          , and_dcpl_367 , and_dcpl_370 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1
          <= 6'b000000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_4_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[6]),
          (operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6[0]), (z_out_36[6]), {and_dcpl_243
          , and_dcpl_373 , and_dcpl_376 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1
          <= MUX1HOT_v_6_4_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[5:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[5:0]),
          ({operator_ac_float_cctor_m_9_lpi_1_dfm_1_5_4 , operator_ac_float_cctor_m_9_lpi_1_dfm_1_3_0}),
          (z_out_36[5:0]), {and_dcpl_243 , and_dcpl_373 , and_dcpl_376 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_5_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_0
          <= MUX1HOT_s_1_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[6]),
          (operator_ac_float_cctor_m_10_lpi_1_dfm_1_10_6[0]), (z_out_37[6]), {and_dcpl_243
          , and_dcpl_399 , and_dcpl_402 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_1
          <= MUX1HOT_v_2_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[5:4]),
          operator_ac_float_cctor_m_10_lpi_1_dfm_1_5_4, (z_out_37[5:4]), {and_dcpl_243
          , and_dcpl_399 , and_dcpl_402 , and_dcpl_192});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2
          <= MUX1HOT_v_4_4_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_6_sva_1[3:0]),
          operator_ac_float_cctor_m_10_lpi_1_dfm_1_3_0, (z_out_37[3:0]), {and_dcpl_243
          , and_dcpl_399 , and_dcpl_402 , and_dcpl_192});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_or_7_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0 <= MUX_s_1_2_2(and_1755_nl,
          (z_out_70[4]), and_dcpl_194);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1 <= MUX_v_4_2_2(nor_571_nl,
          (z_out_70[3:0]), and_dcpl_194);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_1_or_8_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0 <= MUX_s_1_2_2(and_1757_nl,
          (z_out_68[4]), and_dcpl_194);
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1 <= MUX_v_4_2_2(nor_569_nl,
          (z_out_68[3:0]), and_dcpl_194);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_6_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_6_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6]),
          (operator_ac_float_cctor_m_7_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[6]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          (z_out_38[6]), (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_254 , and_dcpl_257 , and_dcpl_199 , and_dcpl_194
          , and_dcpl_215});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1
          <= MUX1HOT_v_2_6_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[5:4]),
          operator_ac_float_cctor_m_7_lpi_1_dfm_1_5_4, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[5:4]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          (z_out_38[5:4]), (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:4]),
          {and_dcpl_243 , and_dcpl_254 , and_dcpl_257 , and_dcpl_199 , and_dcpl_194
          , and_dcpl_215});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2
          <= MUX1HOT_v_4_6_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[3:0]),
          operator_ac_float_cctor_m_7_lpi_1_dfm_1_3_0, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_3_sva_1[3:0]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          (z_out_38[3:0]), (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          {and_dcpl_243 , and_dcpl_254 , and_dcpl_257 , and_dcpl_199 , and_dcpl_194
          , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
          <= 6'b000000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_7_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_6_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[6]),
          (operator_ac_float_cctor_m_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[6]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          (z_out_35[6]), (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_361 , and_dcpl_364 , and_dcpl_199 , and_dcpl_194
          , and_dcpl_215});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1
          <= MUX1HOT_v_6_6_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_itm[5:0]),
          ({operator_ac_float_cctor_m_lpi_1_dfm_1_5_4 , operator_ac_float_cctor_m_lpi_1_dfm_1_3_0}),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_sva_1[5:0]),
          (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:0]),
          (z_out_35[5:0]), (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:0]),
          {and_dcpl_243 , and_dcpl_361 , and_dcpl_364 , and_dcpl_199 , and_dcpl_194
          , and_dcpl_215});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
          <= 6'b000000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_8_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_5_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6]),
          (operator_ac_float_cctor_m_9_lpi_1_dfm_1_10_6[0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[6]),
          (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_373 , and_dcpl_376 , and_dcpl_199 , and_dcpl_194});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1
          <= MUX1HOT_v_6_5_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[5:0]),
          ({operator_ac_float_cctor_m_9_lpi_1_dfm_1_5_4 , operator_ac_float_cctor_m_9_lpi_1_dfm_1_3_0}),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_5_sva_1[5:0]),
          (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:0]),
          (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:0]),
          {and_dcpl_243 , and_dcpl_373 , and_dcpl_376 , and_dcpl_199 , and_dcpl_194});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
          <= 1'b0;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
          <= 2'b00;
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2
          <= 4'b0000;
    end
    else if ( ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_and_9_ssc
        ) begin
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_0
          <= MUX1HOT_s_1_5_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[6]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[6]),
          (operator_ac_float_cctor_m_12_lpi_1_dfm_1_10_6[0]), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[6]),
          (MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[6]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_192 , and_dcpl_195});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_1
          <= MUX1HOT_v_2_5_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[5:4]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[5:4]),
          operator_ac_float_cctor_m_12_lpi_1_dfm_1_5_4, (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[5:4]),
          (MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[5:4]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_192 , and_dcpl_195});
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2
          <= MUX1HOT_v_4_5_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_itm[3:0]),
          (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op2_m_8_sva_1[3:0]),
          operator_ac_float_cctor_m_12_lpi_1_dfm_1_3_0, (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_acc_itm[3:0]),
          (MAC_1_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          {and_dcpl_243 , and_dcpl_392 , and_dcpl_395 , and_dcpl_192 , and_dcpl_195});
    end
  end
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl
      = ~((MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_itm[12]) | i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl = (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_3_lshift_itm[12])
      & (~ i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_nor_15_nl
      = ~((MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_itm[12]) | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_and_31_nl = (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_2_lshift_itm[12])
      & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_unequal_tmp_16);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_6_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_l_qif_mux_7_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_4_else_r_ac_float_4_else_r_ac_float_4_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_6_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_3_else_r_ac_float_3_else_r_ac_float_3_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_l_qif_mux_7_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_2_else_r_ac_float_2_else_r_ac_float_2_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_1_else_r_ac_float_1_else_r_ac_float_1_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl =
      MUX_s_1_2_2((MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_2_nl =
      MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[0]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[1]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_2_nl &
      (~ MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_13_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_13_nl &
      (~ MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl = MUX_s_1_2_2((MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl = MUX_s_1_2_2((MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl = MUX_s_1_2_2((MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl = MUX_s_1_2_2((MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl = MUX_s_1_2_2((MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl = MUX_s_1_2_2((MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl = MUX_s_1_2_2((MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl = MUX_s_1_2_2((MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl = MUX_s_1_2_2((MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl = MUX_s_1_2_2((MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl = MUX_s_1_2_2((MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl = MUX_s_1_2_2((MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl = MUX_s_1_2_2((MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl = MUX_s_1_2_2((MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb;
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl = MUX_s_1_2_2((MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl
      = result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl & result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb;
  assign and_1233_nl = nor_98_cse & (~((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      | MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1236_nl = nor_98_cse & (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1239_nl = (~ (fsm_output[2])) & (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_nl = (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_209 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_24_nl = (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_209 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_25_nl = (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[1]))
      & and_dcpl_199 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_26_nl = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[1])
      & and_dcpl_199 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_27_nl = (~ (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_192 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_28_nl = (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_192 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_29_nl = (~ (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1425 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_30_nl = (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1425 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_31_nl = (~ (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1427 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_32_nl = (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1427 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_33_nl = (~ (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1428 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_34_nl = (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1428 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_35_nl = (~ (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1429 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_36_nl = (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1429 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_37_nl = (~ (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1430 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_38_nl = (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1430 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_39_nl = (~ (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1431 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_40_nl = (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1431 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_41_nl = (~ (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1432 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_42_nl = (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1432 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_43_nl = (~ (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1433 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_44_nl = (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1433 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_45_nl = (~ (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1434 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_46_nl = (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1434 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_47_nl = (~ (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1435 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_48_nl = (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1435 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_49_nl = (~ (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1436 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_50_nl = (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1436 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_51_nl = (~ (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1437 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_52_nl = (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1437 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_53_nl = (~ (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1438 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_54_nl = (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1438 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_55_nl = (~ (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1439 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_56_nl = (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1439 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_57_nl = (~ (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1440 & (~ or_1011_tmp);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_58_nl = (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1440 & (~ or_1011_tmp);
  assign mux1h_12_nl = MUX1HOT_v_4_42_2((MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[3:0]), (z_out_4[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_115,
      leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_127, (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0, (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_2_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_3_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_4_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_5_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_6_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_7_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_8_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_9_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_10_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_11_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_12_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_13_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_14_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_15_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_16_result_imag_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      {and_dcpl_186 , and_1233_nl , and_1236_nl , and_1239_nl , and_dcpl_194 , and_dcpl_195
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_24_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_25_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_26_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_27_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_28_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_29_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_30_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_31_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_32_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_33_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_34_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_35_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_36_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_37_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_38_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_39_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_40_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_41_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_42_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_43_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_44_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_45_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_46_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_47_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_48_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_49_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_50_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_51_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_52_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_53_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_54_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_55_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_56_nl
      , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_57_nl , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_and_58_nl});
  assign not_1835_nl = ~ or_1011_tmp;
  assign and_1033_nl = and_dcpl_937 & nor_98_cse & (~((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      | MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_1036_nl = and_dcpl_937 & nor_98_cse & (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  assign and_1039_nl = and_dcpl_188 & (~ (fsm_output[2])) & (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      & (~ mux_123_itm);
  assign and_951_nl = and_dcpl_937 & nor_98_cse & (~((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      | MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_954_nl = and_dcpl_937 & nor_98_cse & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1;
  assign and_957_nl = and_dcpl_188 & (~ (fsm_output[2])) & (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      & (~ mux_123_itm);
  assign mux_350_nl = MUX_s_1_2_2(or_tmp_111, or_tmp_107, fsm_output[0]);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, or_tmp_102, fsm_output[3]);
  assign mux_352_nl = MUX_s_1_2_2(mux_tmp_121, mux_351_nl, fsm_output[2]);
  assign and_972_nl = nor_98_cse & (~((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_975_nl = nor_98_cse & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_978_nl = (~ (fsm_output[2])) & (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign and_1043_nl = nor_98_cse & (~((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1046_nl = nor_98_cse & (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1049_nl = (~ (fsm_output[2])) & (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign and_1150_nl = nor_98_cse & (~((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1153_nl = nor_98_cse & (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1156_nl = (~ (fsm_output[2])) & (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign and_1198_nl = nor_98_cse & (~((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1201_nl = nor_98_cse & (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1204_nl = (~ (fsm_output[2])) & (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign and_1243_nl = nor_98_cse & (~((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1246_nl = nor_98_cse & (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1249_nl = (~ (fsm_output[2])) & (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_9_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[54:50]);
  assign MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign and_1782_nl = and_dcpl_194 & nor_559_m1c;
  assign and_1783_nl = and_dcpl_195 & nor_559_m1c;
  assign and_1784_nl = and_dcpl_198 & nor_559_m1c;
  assign or_nl = ((~ MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1)
      & and_1785_m1c) | or_dcpl_543;
  assign and_2626_nl = MAC_2_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_1_itm_6_1
      & and_1785_m1c;
  assign mux1h_8_nl = MUX1HOT_v_6_8_2(MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp,
      (z_out_12[5:0]), z_out_6, (z_out_9[5:0]), 6'b110000, MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_else_1_qelse_acc_itm,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6, {and_dcpl_186
      , and_dcpl_209 , and_1782_nl , and_1783_nl , and_1784_nl , or_nl , and_2626_nl
      , and_dcpl_213});
  assign not_1826_nl = ~ or_dcpl_544;
  assign and_1779_nl = MUX_v_6_2_2(6'b000000, mux1h_8_nl, not_1826_nl);
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_10_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign or_1074_nl = (and_dcpl_194 & nor_560_m1c) | (and_dcpl_212 & nor_560_m1c);
  assign or_1075_nl = (and_dcpl_195 & nor_560_m1c) | (and_dcpl_198 & nor_560_m1c);
  assign mux1h_9_nl = MUX1HOT_v_6_6_2(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
      MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      z_out_6, (z_out_15[5:0]), r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_qr_5_0_3_lpi_1_dfm_mx0w6,
      6'b110000, {and_dcpl_186 , and_dcpl_209 , or_1074_nl , or_1075_nl , and_dcpl_213
      , or_dcpl_546});
  assign not_1825_nl = ~ or_dcpl_548;
  assign and_1771_nl = MUX_v_6_2_2(6'b000000, mux1h_9_nl, not_1825_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_7_nl = MUX_v_2_2_2((z_out_27[6:5]),
      (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl
      = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_7_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl
      = MUX_v_2_2_2(2'b00, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_seb);
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_2_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_2_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_10_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_10_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_72 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_88 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_98 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[0])));
  assign or_897_nl = MAC_2_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp
      | MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp;
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_10_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_10_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_71 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_86 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_96 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_if_nand_1_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_104 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])));
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_15_nl =
      MUX_s_1_2_2((MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_15_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_15_nl & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_14_nl
      = MUX_s_1_2_2((MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_14_nl &
      (~ MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl = MUX_s_1_2_2((MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl = MUX_s_1_2_2((MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_1_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_1_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl = MUX_s_1_2_2((MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_2_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_2_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_2_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl = MUX_s_1_2_2((MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_3_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_3_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_3_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl = MUX_s_1_2_2((MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_4_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_4_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_4_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl = MUX_s_1_2_2((MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_5_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_5_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_5_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl = MUX_s_1_2_2((MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_6_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_6_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_6_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl = MUX_s_1_2_2((MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_7_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_7_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_7_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl = MUX_s_1_2_2((MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_8_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_8_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_8_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl = MUX_s_1_2_2((MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_9_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_9_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_9_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl = MUX_s_1_2_2((MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_10_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_10_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_10_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl = MUX_s_1_2_2((MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_11_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_11_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_11_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl = MUX_s_1_2_2((MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_12_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_12_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_12_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl = MUX_s_1_2_2((MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_13_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_13_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_13_seb;
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl = MUX_s_1_2_2((MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_14_nl
      = result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_14_nl & result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_14_seb;
  assign and_960_nl = nor_98_cse & (~((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2])
      | MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_963_nl = nor_98_cse & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_966_nl = (~ (fsm_output[2])) & (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_nl = (~ (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_209 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl = (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_209 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_3_nl = (~ (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_192 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl = (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_192 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_5_nl = (~ (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1425 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_6_nl = (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1425 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl = (~ (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1427 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl = (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1427 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_9_nl = (~ (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1428 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_10_nl = (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1428 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_nl = (~ (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1429 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_12_nl = (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1429 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl = (~ (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1430 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl = (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1430 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl = (~ (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1431 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_16_nl = (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1431 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_17_nl = (~ (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1432 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_18_nl = (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1432 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_19_nl = (~ (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1433 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_20_nl = (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1433 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_21_nl = (~ (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1434 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_22_nl = (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1434 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl = (~ (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1435 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_24_nl = (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1435 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_25_nl = (~ (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1436 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_26_nl = (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1436 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_27_nl = (~ (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1437 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_28_nl = (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1437 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_29_nl = (~ (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1438 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_30_nl = (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1438 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_31_nl = (~ (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1439 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_32_nl = (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1439 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_33_nl = (~ (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1440 & (~ or_1065_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_34_nl = (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1440 & (~ or_1065_tmp);
  assign mux1h_13_nl = MUX1HOT_v_4_40_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg[3:0]), (z_out_2[3:0]), leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_113,
      leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_126, (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_mx0w2_3_0,
      (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_2_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_3_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_4_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_5_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_6_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_7_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_8_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_9_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_10_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_11_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_12_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_13_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_14_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_15_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_16_result_real_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      {and_960_nl , and_963_nl , and_966_nl , and_dcpl_194 , and_dcpl_195 , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_2_nl , and_dcpl_199
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_3_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_5_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_6_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_9_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_10_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_11_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_12_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_13_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_16_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_17_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_18_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_19_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_20_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_21_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_22_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_24_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_25_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_26_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_27_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_28_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_29_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_30_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_31_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_32_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_33_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_34_nl});
  assign not_1837_nl = ~ or_1065_tmp;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl = (~ nor_474_tmp)
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl = nor_474_tmp
      & and_dcpl_209;
  assign nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_4_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[29:25]);
  assign MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_9_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[54:50]);
  assign MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_11_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign mux_110_nl = MUX_s_1_2_2(or_tmp_104, or_tmp_102, fsm_output[3]);
  assign mux_108_nl = MUX_s_1_2_2(mux_tmp_101, or_dcpl_196, fsm_output[0]);
  assign mux_109_nl = MUX_s_1_2_2(mux_108_nl, or_tmp_102, fsm_output[3]);
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_10_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign and_1832_nl = and_dcpl_195 & nor_551_m1c;
  assign and_1833_nl = and_dcpl_198 & nor_551_m1c;
  assign mux1h_nl = MUX1HOT_v_6_6_2(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
      MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1, (z_out_9[5:0]),
      z_out_6, 6'b110000, {and_dcpl_186 , and_dcpl_209 , and_dcpl_199 , and_1832_nl
      , and_1833_nl , or_dcpl_526});
  assign not_1834_nl = ~ or_dcpl_527;
  assign and_1827_nl = MUX_v_6_2_2(6'b000000, mux1h_nl, not_1834_nl);
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_11_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign and_1825_nl = and_dcpl_195 & nor_552_m1c;
  assign and_1826_nl = and_dcpl_198 & nor_552_m1c;
  assign mux1h_1_nl = MUX1HOT_v_6_6_2(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
      MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1, (z_out_11[5:0]),
      (z_out_5[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_209 , and_dcpl_199 , and_1825_nl
      , and_1826_nl , or_dcpl_528});
  assign not_1833_nl = ~ or_dcpl_529;
  assign and_1820_nl = MUX_v_6_2_2(6'b000000, mux1h_1_nl, not_1833_nl);
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_11_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign and_1818_nl = and_dcpl_195 & nor_553_m1c;
  assign and_1819_nl = and_dcpl_198 & nor_553_m1c;
  assign mux1h_2_nl = MUX1HOT_v_6_6_2(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w2, (z_out_12[5:0]),
      (z_out_11[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_209 , and_dcpl_199 , and_1818_nl
      , and_1819_nl , or_dcpl_530});
  assign not_1832_nl = ~ or_dcpl_531;
  assign and_1813_nl = MUX_v_6_2_2(6'b000000, mux1h_2_nl, not_1832_nl);
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_13_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign and_1811_nl = and_dcpl_195 & nor_554_m1c;
  assign and_1812_nl = and_dcpl_198 & nor_554_m1c;
  assign mux1h_3_nl = MUX1HOT_v_6_5_2(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
      z_out_3, (z_out_20[5:0]), (z_out_16[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_199
      , and_1811_nl , and_1812_nl , or_dcpl_532});
  assign not_1831_nl = ~ or_dcpl_533;
  assign and_1807_nl = MUX_v_6_2_2(6'b000000, mux1h_3_nl, not_1831_nl);
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_13_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign and_1805_nl = and_dcpl_195 & nor_555_m1c;
  assign and_1806_nl = and_dcpl_198 & nor_555_m1c;
  assign mux1h_4_nl = MUX1HOT_v_6_5_2(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1, (z_out_4[5:0]),
      (z_out_21[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_199 , and_1805_nl , and_1806_nl
      , or_dcpl_534});
  assign not_1830_nl = ~ or_dcpl_535;
  assign and_1801_nl = MUX_v_6_2_2(6'b000000, mux1h_4_nl, not_1830_nl);
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_11_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign and_1793_nl = and_dcpl_195 & nor_557_m1c;
  assign and_1794_nl = and_dcpl_198 & nor_557_m1c;
  assign mux1h_6_nl = MUX1HOT_v_6_4_2(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
      (z_out_18[5:0]), (z_out_4[5:0]), 6'b110000, {and_dcpl_186 , and_1793_nl , and_1794_nl
      , or_dcpl_538});
  assign not_1828_nl = ~ or_dcpl_539;
  assign and_1791_nl = MUX_v_6_2_2(6'b000000, mux1h_6_nl, not_1828_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_37_nl =
      (~ nor_489_tmp) & and_dcpl_209;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_38_nl =
      nor_489_tmp & and_dcpl_209;
  assign and_1135_nl = nor_98_cse & (~((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      | MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_260;
  assign and_1138_nl = nor_98_cse & (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_260;
  assign and_1141_nl = (~ (fsm_output[2])) & (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_260;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_1_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_1_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_1_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_2_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_2_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_2_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_2_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_2_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_2_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_2_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_3_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_3_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_3_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_3_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_3_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_3_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_3_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_4_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_4_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_4_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_4_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_4_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_4_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_5_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_5_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_5_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_5_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_5_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_5_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_6_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_6_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_6_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_6_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_6_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_6_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_7_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_7_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_7_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_7_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_7_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_7_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_8_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_actual_max_shift_left_acc_psp_8_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_8_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_psp_8_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_acc_psp_8_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_15_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_15_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_15_sva_1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_sva_mx0w1[6:4])
      + 3'b001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      = ~((~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_nl
      = MUX1HOT_v_5_3_2((z_out_27[4:0]), 5'b10000, (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_16_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_seb);
  assign nand_54_nl = ~(or_972_cse & (fsm_output[1:0]==2'b11));
  assign or_744_nl = (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5:4]!=2'b01)
      | (fsm_output[0]))) | (fsm_output[1]);
  assign mux_481_nl = MUX_s_1_2_2(nand_54_nl, or_744_nl, fsm_output[3]);
  assign or_741_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5:4]!=2'b00)
      | (fsm_output[1:0]!=2'b00);
  assign nor_71_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm));
  assign mux_480_nl = MUX_s_1_2_2(or_tmp_20, or_741_nl, nor_71_nl);
  assign or_742_nl = (fsm_output[3]) | mux_480_nl;
  assign mux_482_nl = MUX_s_1_2_2(mux_481_nl, or_742_nl, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl = (mux_482_nl
      | or_dcpl_207) & and_362_ssc;
  assign and_1469_nl = or_972_cse & and_dcpl_976 & and_362_ssc;
  assign and_1472_nl = (and_dcpl_1463 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_14_itm)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0)
      & and_dcpl_1054 & and_362_ssc;
  assign and_1473_nl = and_dcpl_1366 & and_dcpl_985;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_1_nl =
      MUX1HOT_s_1_4_2((MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[4]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_1[0]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[4]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_1_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_3_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c3});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_28_nl =
      MUX1HOT_v_4_4_2((MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[3:0]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_12_sva_rsp_1_rsp_2,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[3:0]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_1_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_3_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_mx0c3});
  assign nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_9_nl = ((~
      or_982_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c1)
      | ((~ or_981_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c2)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c7;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_5_nl = or_982_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_7_nl = or_981_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva_mx0c2;
  assign nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_5_nl =
      MUX1HOT_s_1_23_2((MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0[4]),
      (operator_ac_float_cctor_e_62_lpi_1_dfm[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0[4]),
      (operator_ac_float_cctor_e_64_lpi_1_dfm[4]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva[4]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva[4]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_4, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva[4]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[4]), operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[4]), {and_dcpl_189
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_9_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_11_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c3
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_13_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c7
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c10
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c11
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c12
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c13
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c14
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c15
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c16
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c17
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c18
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c19
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c20
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c21
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c22
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c23});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_18_nl =
      MUX1HOT_v_4_23_2((MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_3_lpi_1_dfm_1_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_3_lpi_1_dfm_1_5_0[3:0]),
      (operator_ac_float_cctor_e_62_lpi_1_dfm[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_12_lpi_1_dfm_1_5_0[3:0]),
      (operator_ac_float_cctor_e_64_lpi_1_dfm[3:0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_9_sva_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0,
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1, operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[3:0]), operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[3:0]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_9_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_11_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c3
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_13_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c7
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_14_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c10
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c11
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c12
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c13
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c14
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c15
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c16
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c17
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c18
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c19
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c20
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c21
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c22
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_11_sva_mx0c23});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_11_nl = ((~
      or_980_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c1)
      | ((~ or_979_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c2)
      | ((~ or_994_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c3)
      | ((~ or_993_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c4)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c8;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_17_nl = or_980_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_19_nl = or_979_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_21_nl = or_994_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c3;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_23_nl = or_993_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_12_sva_mx0c4;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl = MUX_s_1_2_2((MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_mux_nl & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_4 &
      (~ MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_15_nl
      = MUX_s_1_2_2((MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_15_nl &
      (~ MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_3_nl =
      MUX1HOT_s_1_5_2((MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[4]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_and_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_4_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_15_nl,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[4]),
      {and_dcpl_189 , and_dcpl_209 , and_dcpl_199 , and_dcpl_192 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c5});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_14_nl = (~
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_15_nl = (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_16_nl = (~
      (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]))
      & and_dcpl_192;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_17_nl = (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      & and_dcpl_192;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_4_nl =
      MUX1HOT_v_4_8_2((MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[3:0]), (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_23_3_0, (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_110, (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[3:0]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_15_nl , and_dcpl_199
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_16_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_17_nl
      , and_dcpl_194 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c5});
  assign nor_566_nl = ~(MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_4_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_mx0c6));
  assign or_1068_nl = (and_dcpl_209 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_nor_1_seb))
      | (MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs &
      and_dcpl_192) | (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs
      & and_dcpl_199);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_12_nl = ((~
      or_978_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c1)
      | ((~ or_977_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c2)
      | ((~ or_992_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c4)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c8;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_25_nl = or_978_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_27_nl = or_977_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_29_nl = or_992_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_13_sva_mx0c4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_11_nl =
      MUX1HOT_s_1_8_2((MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0[4]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0[4]),
      (operator_ac_float_cctor_e_34_lpi_1_dfm[4]), (operator_ac_float_cctor_e_19_lpi_1_dfm[4]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0[0]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_31_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_33_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c3
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_35_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c7});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_mux1h_29_nl =
      MUX1HOT_v_4_8_2((MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_7_lpi_1_dfm_1_5_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_7_lpi_1_dfm_1_5_0[3:0]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1_5_0[3:0]),
      (operator_ac_float_cctor_e_34_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_19_lpi_1_dfm[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_31_ssc
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_33_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c3
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_35_ssc , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_mx0c7});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_or_14_nl = ((~
      or_974_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c1)
      | ((~ or_973_cse) & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c2)
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c6;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_37_nl = or_974_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_and_39_nl = or_973_cse
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_15_sva_mx0c2;
  assign nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_11_sva[21]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_9_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_10_sva[21]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_11_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl = ~((operator_ac_float_cctor_m_31_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_7_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_8_sva[21]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_8_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_9_sva[21]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_16_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_3_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_13_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl = ~((operator_ac_float_cctor_m_33_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_14_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl = ~((operator_ac_float_cctor_m_34_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_11_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_61_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign MAC_12_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_nl = ~((operator_ac_float_cctor_m_32_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_1_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_2_sva[21]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign MAC_12_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_62_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_2_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_3_sva[21]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign MAC_13_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_63_lpi_1_dfm_mx0w0!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_3_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_4_sva[21]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign MAC_14_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_64_lpi_1_dfm_mx0w0!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_4_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_r_m_5_sva[21]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nor_itm);
  assign MAC_15_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_nl = ~((operator_ac_float_cctor_m_65_lpi_1_dfm_mx0w0!=11'b00000000000));
  assign MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_3_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_3_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_11_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | ac_float_cctor_operator_return_59_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_70 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_sva_0));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_84 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_4_sva_3_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_94 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2[0])));
  assign or_899_nl = MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_3_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | ac_float_cctor_operator_return_29_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_73 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_82 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_3_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_92 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1[0])));
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_4_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_4_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_12_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | ac_float_cctor_operator_return_60_sva;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_80 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_6_sva_3_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_14_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_91 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1[0])));
  assign MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_4_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | ac_float_cctor_operator_return_30_sva;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_78 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_3_0[0])));
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_15_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_90 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_1_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_2_sva[21]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_5_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_5_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = ac_float_cctor_operator_return_46_sva_mx0w2
      | ac_float_cctor_operator_return_61_sva;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_76 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_10_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_11_sva[21]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_5_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = ac_float_cctor_operator_return_16_sva_mx0w2
      | ac_float_cctor_operator_return_31_sva;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_74 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_10_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_99 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_11_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_12_sva[21]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_6_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_6_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = ac_float_cctor_operator_return_47_sva_mx0w2
      | ac_float_cctor_operator_return_62_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_5_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_81 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_12_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_13_sva[21]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_6_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = ac_float_cctor_operator_return_17_sva_mx0w2
      | ac_float_cctor_operator_return_32_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_1_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_89 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_11_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_97 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_13_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_14_sva[21]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = MAC_7_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp
      | MAC_7_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp;
  assign MAC_15_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = ac_float_cctor_operator_return_48_sva_mx0w2
      | ac_float_cctor_operator_return_63_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_2_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_87 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_4_sva[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_12_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_95 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_14_sva_0));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_2_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_3_sva[21]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_7_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = ac_float_cctor_operator_return_2_sva_mx0w2
      | ac_float_cctor_operator_return_3_sva;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_3_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_85 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_5_sva[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_13_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_93 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_15_sva_0));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_3_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_4_sva[21]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign or_898_nl = MAC_8_ac_float_cctor_operator_3_ac_float_cctor_operator_3_nor_tmp
      | MAC_8_ac_float_cctor_operator_2_ac_float_cctor_operator_2_nor_tmp;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_4_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_83 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_6_sva[0])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_9_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_101 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva[0])));
  assign MAC_6_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl
      = ~((operator_r_m_6_lpi_1_dfm_mx0w5_10_6!=5'b00000) | (operator_r_m_6_lpi_1_dfm_mx0w5_5_4!=2'b00)
      | (operator_r_m_6_lpi_1_dfm_mx0w5_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_4_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_5_sva[21]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp
      | MAC_8_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_6_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_79 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_8_sva[0])));
  assign MAC_7_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl
      = ~((operator_r_m_7_lpi_1_dfm_mx0w4_10_6!=5'b00000) | (operator_r_m_7_lpi_1_dfm_mx0w4_5_4!=2'b00)
      | (operator_r_m_7_lpi_1_dfm_mx0w4_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_5_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_6_sva[21]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_nl = ac_float_cctor_operator_return_42_sva_mx0w1
      | ac_float_cctor_operator_return_57_sva_mx0w1;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_7_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_77 & (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva[0])));
  assign MAC_8_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl
      = ~((operator_r_m_8_lpi_1_dfm_mx0w6_10_6!=5'b00000) | (operator_r_m_8_lpi_1_dfm_mx0w6_5_4!=2'b00)
      | (operator_r_m_8_lpi_1_dfm_mx0w6_3_0!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nand_6_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_r_m_7_sva[21]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_if_nor_itm);
  assign MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_nl = ac_float_cctor_operator_return_12_sva_mx0w1
      | ac_float_cctor_operator_return_27_sva_mx0w1;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_8_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_75 & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_10_sva_0));
  assign MAC_9_my_complex_float_t_cctor_real_operator_my_complex_float_t_cctor_real_operator_nor_nl
      = ~((operator_r_m_9_lpi_1_dfm_mx0w6_10_6!=5'b00000) | (operator_r_m_9_lpi_1_dfm_mx0w6_5_4!=2'b00)
      | (operator_r_m_9_lpi_1_dfm_mx0w6_3_0!=4'b0000));
  assign nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_38_nl = ~ MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_7_nl
      = MUX_v_5_2_2(5'b00000, z_out_31, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_38_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_16_nl = or_487_rgt & (~ and_dcpl_192);
  assign mux_442_nl = MUX_s_1_2_2(not_tmp_307, mux_tmp_150, fsm_output[3]);
  assign mux_443_nl = MUX_s_1_2_2(mux_442_nl, mux_tmp_149, fsm_output[2]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_8_nl =
      MUX_s_1_2_2((MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl
      = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_8_nl &
      (~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_6_nl
      = MUX1HOT_s_1_5_2((MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[4]), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_8_nl,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0[0]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_mx0w1[4]), {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , and_1331_rgt , and_dcpl_192});
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_36_nl
      = MUX_v_4_2_2((MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_82_nl = ~ MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl
      = MUX_v_4_2_2(4'b0000, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_36_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_not_82_nl);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_operator_13_2_true_AC_TRN_AC_WRAP_1_mux1h_13_nl
      = MUX1HOT_v_4_5_2((MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[3:0]), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_23_nl,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_mx0w1[3:0]), {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , and_1331_rgt , and_dcpl_192});
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_8_sva_mx0w1[5:4]) + 2'b01;
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_7_sva_mx0w1[5:4]) + 2'b01;
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_6_sva_mx0w1[5:4]) + 2'b01;
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_5_sva_mx0w1[5:4]) + 2'b01;
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1[5:4]) + 2'b01;
  assign nl_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_3_sva_mx0w1[5:4]) + 2'b01;
  assign nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl
      = (z_out[5:4]) + 2'b01;
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl
      = nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (z_out_29[5:4]) + 2'b01;
  assign MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_16_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (z_out_30[5:4]) + 2'b01;
  assign MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_15_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (z_out_28[5:4]) + 2'b01;
  assign MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:4]) + 2'b01;
  assign MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl
      = (z_out_1[5:4]) + 2'b01;
  assign MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl
      = nl_MAC_1_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_nl[1:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_1_nl =
      MUX1HOT_s_1_8_2((MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[4]), (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[4]), (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[4]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[4]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_2_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_3_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_4_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_5_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_6_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_7_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c5});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_5_nl =
      MUX1HOT_v_4_9_2((MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[3:0]), (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3:0]), (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_2_sva_4_0[3:0]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[3:0]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_sdt[3:0]),
      leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_112, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]),
      {and_dcpl_189 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_2_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_3_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_4_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_5_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_6_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_and_7_cse , and_dcpl_194
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c5});
  assign nor_574_nl = ~(MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_mux1h_5_nl,
      4'b1111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_mx0c6));
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_11_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign mux_125_nl = MUX_s_1_2_2(or_tmp_111, or_dcpl_207, fsm_output[0]);
  assign mux_126_nl = MUX_s_1_2_2(mux_125_nl, or_tmp_102, fsm_output[3]);
  assign mux_128_nl = MUX_s_1_2_2(mux_tmp_121, mux_126_nl, fsm_output[2]);
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_12_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_13_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_14_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_13_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign nor_218_nl = ~((~ (fsm_output[3])) | (fsm_output[0]) | (fsm_output[1]));
  assign nor_219_nl = ~((fsm_output[3]) | mux_tmp_31);
  assign mux_130_nl = MUX_s_1_2_2(nor_218_nl, nor_219_nl, fsm_output[2]);
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_12_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_12_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_12_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(input_real_e_rsci_idat)
      + conv_s2s_5_6(taps_real_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_0_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[9:5]);
  assign MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_0_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[9:5]);
  assign MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_14_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign and_1799_nl = and_dcpl_195 & nor_556_m1c;
  assign and_1800_nl = and_dcpl_198 & nor_556_m1c;
  assign mux1h_5_nl = MUX1HOT_v_6_5_2(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl,
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_4_sva_mx0w1, (z_out_16[5:0]),
      (z_out_25[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_192 , and_1799_nl , and_1800_nl
      , or_dcpl_536});
  assign not_1829_nl = ~ or_dcpl_537;
  assign and_1795_nl = MUX_v_6_2_2(6'b000000, mux1h_5_nl, not_1829_nl);
  assign or_337_nl = (fsm_output[3]) | nor_137_cse;
  assign mux_148_nl = MUX_s_1_2_2(or_tmp_20, or_337_nl, fsm_output[2]);
  assign and_236_nl = (~ mux_148_nl) & and_dcpl_206;
  assign mux_551_nl = MUX_s_1_2_2(mux_536_cse, or_dcpl_200, fsm_output[2]);
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_14_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl = MUX_v_6_2_2(6'b110000,
      (z_out_8[5:0]), MAC_6_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_20_nl
      = MUX_v_6_2_2(6'b000000, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_16_nl,
      MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(input_imag_e_rsci_idat)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl = MUX_v_6_2_2(6'b110000,
      (z_out_10[5:0]), MAC_7_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_21_nl
      = MUX_v_6_2_2(6'b000000, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_19_nl,
      MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(input_real_e_rsci_idat)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl = MUX_v_6_2_2(6'b110000,
      (z_out_7[5:0]), MAC_8_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_22_nl
      = MUX_v_6_2_2(6'b000000, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_nl,
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs);
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(input_imag_e_rsci_idat)
      + conv_s2s_5_6(taps_real_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl = MUX_v_6_2_2(6'b110000,
      (z_out_25[5:0]), MAC_9_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_23_nl
      = MUX_v_6_2_2(6'b000000, r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_nl,
      MAC_9_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_or_svs);
  assign nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_0_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[9:5]);
  assign MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_7_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = (~ (MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl
      = nl_MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_qif_acc_nl[4:0];
  assign nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = nl_MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_33_nl =
      or_736_rgt & ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_mx0c2;
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_nl = MUX1HOT_s_1_19_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0[4]),
      (operator_ac_float_cctor_e_61_lpi_1_dfm[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0[4]),
      (operator_ac_float_cctor_e_63_lpi_1_dfm[4]), (operator_ac_float_cctor_e_31_lpi_1_dfm[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[4]),
      (operator_ac_float_cctor_e_62_lpi_1_dfm[4]), (operator_ac_float_cctor_e_64_lpi_1_dfm[4]),
      (operator_ac_float_cctor_e_65_lpi_1_dfm[4]), (operator_ac_float_cctor_e_14_lpi_1_dfm[4]),
      (operator_ac_float_cctor_e_19_lpi_1_dfm[4]), (operator_ac_float_cctor_e_29_lpi_1_dfm[4]),
      (operator_ac_float_cctor_e_3_lpi_1_dfm[4]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[4]),
      (operator_ac_float_cctor_e_33_lpi_1_dfm[4]), (operator_ac_float_cctor_e_34_lpi_1_dfm[4]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0,
      {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_3_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_5_itm
      , and_1488_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_7_itm
      , and_1494_itm , and_1496_itm , and_1499_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_itm
      , and_1504_itm , and_1507_itm , and_1510_itm , and_1513_itm , and_1516_itm
      , and_1519_itm , and_1522_itm , and_1525_itm , and_1528_itm , and_1531_itm
      , and_1534_itm});
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_8_nl = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_nl
      & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_itm);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_1_nl =
      MUX1HOT_v_4_19_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_qr_6_0_2_lpi_1_dfm_1_5_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_2_lpi_1_dfm_1_5_0[3:0]),
      (operator_ac_float_cctor_e_61_lpi_1_dfm[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_qr_6_0_11_lpi_1_dfm_1_5_0[3:0]),
      (operator_ac_float_cctor_e_63_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_31_lpi_1_dfm[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[3:0]),
      (operator_ac_float_cctor_e_62_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_64_lpi_1_dfm[3:0]),
      (operator_ac_float_cctor_e_65_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_14_lpi_1_dfm[3:0]),
      (operator_ac_float_cctor_e_19_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_29_lpi_1_dfm[3:0]),
      (operator_ac_float_cctor_e_3_lpi_1_dfm[3:0]), (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]),
      (operator_ac_float_cctor_e_33_lpi_1_dfm[3:0]), (operator_ac_float_cctor_e_34_lpi_1_dfm[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1,
      {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_3_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_5_itm
      , and_1488_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_7_itm
      , and_1494_itm , and_1496_itm , and_1499_itm , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_and_itm
      , and_1504_itm , and_1507_itm , and_1510_itm , and_1513_itm , and_1516_itm
      , and_1519_itm , and_1522_itm , and_1525_itm , and_1528_itm , and_1531_itm
      , and_1534_itm});
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_1_nl = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_mux1h_1_nl,
      4'b1111, ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_t_or_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl = (~ nor_495_tmp)
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl = nor_495_tmp
      & and_dcpl_209;
  assign or_1097_nl = (((((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5:4]!=2'b00))
      & MAC_16_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) |
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4]))
      & (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | not_tmp_1312;
  assign or_1094_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[4])
      & (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | not_tmp_1312;
  assign mux_552_nl = MUX_s_1_2_2(or_1097_nl, or_1094_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0);
  assign or_1093_nl = (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | not_tmp_1312;
  assign or_1091_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1[2:0]!=3'b000)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0[3:0]!=4'b0000)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0!=2'b00)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1[3]);
  assign mux_553_nl = MUX_s_1_2_2(mux_552_nl, or_1093_nl, or_1091_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl = (~ nor_493_tmp)
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl = nor_493_tmp
      & and_dcpl_209;
  assign or_1108_nl = (((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5:4]!=2'b00))
      & MAC_8_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_or_svs) | (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      | not_tmp_1322;
  assign or_1105_nl = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[4])
      | not_tmp_1322;
  assign mux_554_nl = MUX_s_1_2_2(or_1108_nl, or_1105_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0);
  assign or_1109_nl = (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1[1:0]!=2'b00)
      | (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_0[3:0]!=4'b0000)
      | (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_0!=2'b00)
      | (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_2_sva_10_0_rsp_1_rsp_1[3:2]!=2'b00)
      | mux_554_nl;
  assign mux_555_nl = MUX_s_1_2_2(not_tmp_1322, or_1109_nl, MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_22_nl = (~ nor_487_tmp) & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_23_nl = nor_487_tmp & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_24_nl = (~ nor_485_tmp) & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_25_nl = nor_485_tmp & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_26_nl = (~ nor_519_tmp) & and_dcpl_209;
  assign operator_13_2_true_AC_TRN_AC_WRAP_1_and_27_nl = nor_519_tmp & and_dcpl_209;
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = conv_s2s_5_6(delay_lane_real_e_10_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl[5:0];
  assign or_1076_nl = (and_dcpl_194 & nor_561_m1c) | (and_dcpl_195 & nor_561_m1c);
  assign and_1770_nl = and_dcpl_198 & nor_561_m1c;
  assign mux1h_10_nl = MUX1HOT_v_6_5_2(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_nl,
      MAC_4_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      (z_out_5[5:0]), (z_out_14[5:0]), 6'b110000, {and_dcpl_186 , and_dcpl_209 ,
      or_1076_nl , and_1770_nl , or_dcpl_550});
  assign not_1824_nl = ~ or_dcpl_552;
  assign and_1765_nl = MUX_v_6_2_2(6'b000000, mux1h_10_nl, not_1824_nl);
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = conv_s2s_5_6(delay_lane_imag_e_10_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl[5:0];
  assign and_1762_nl = and_dcpl_194 & nor_562_m1c;
  assign and_1763_nl = and_dcpl_195 & nor_562_m1c;
  assign and_1764_nl = and_dcpl_198 & nor_562_m1c;
  assign mux1h_11_nl = MUX1HOT_v_6_6_2(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_nl,
      MAC_5_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp,
      (z_out_11[5:0]), (z_out_14[5:0]), (z_out_12[5:0]), 6'b110000, {and_dcpl_186
      , and_dcpl_209 , and_1762_nl , and_1763_nl , and_1764_nl , or_dcpl_554});
  assign not_1823_nl = ~ or_dcpl_555;
  assign and_1759_nl = MUX_v_6_2_2(6'b000000, mux1h_11_nl, not_1823_nl);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1[3:0]);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_acc_nl[3:0];
  assign and_1184_nl = nor_98_cse & (~((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      | MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_260;
  assign and_1187_nl = nor_98_cse & (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_260;
  assign and_1190_nl = (~ (fsm_output[2])) & (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_260;
  assign or_1144_nl = (~((~((~(and_dcpl_1554 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_9_itm)))
      | (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])))
      | (~ (fsm_output[2])) | (fsm_output[0]))) | (fsm_output[1]);
  assign nor_787_nl = ~((fsm_output[2:0]!=3'b001));
  assign mux_556_nl = MUX_s_1_2_2(or_1144_nl, nor_787_nl, fsm_output[6]);
  assign nor_788_nl = ~((fsm_output[6]) | (~((~ (fsm_output[2])) | (fsm_output[0])))
      | (fsm_output[1]));
  assign mux_557_nl = MUX_s_1_2_2(mux_556_nl, nor_788_nl, fsm_output[3]);
  assign nor_789_nl = ~((fsm_output[6]) | (~ (fsm_output[0])) | (fsm_output[1]));
  assign nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = conv_s2s_5_6(delay_lane_real_e_4_sva)
      + conv_s2s_5_6(taps_real_e_rsci_idat[29:25]);
  assign MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl = nl_MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_nl[5:0];
  assign or_1126_nl = (fsm_output[1]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      | (~(((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[5:4]!=2'b00))
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_10_itm))));
  assign mux_559_nl = MUX_s_1_2_2(or_1126_nl, (fsm_output[1]), fsm_output[0]);
  assign nor_793_nl = ~((fsm_output[3]) | (~ mux_559_nl));
  assign mux_560_nl = MUX_s_1_2_2(nor_793_nl, nor_794_cse, MAC_11_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign mux_562_nl = MUX_s_1_2_2(mux_561_cse, mux_560_nl, fsm_output[2]);
  assign or_1132_nl = (fsm_output[1]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0
      | (~(((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5:4]!=2'b00))
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_11_itm))));
  assign mux_563_nl = MUX_s_1_2_2(or_1132_nl, (fsm_output[1]), fsm_output[0]);
  assign nor_800_nl = ~((fsm_output[3]) | (~ mux_563_nl));
  assign mux_564_nl = MUX_s_1_2_2(nor_800_nl, nor_794_cse, MAC_12_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5]);
  assign mux_566_nl = MUX_s_1_2_2(mux_561_cse, mux_564_nl, fsm_output[2]);
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = conv_s2s_5_6(delay_lane_imag_e_8_sva)
      + conv_s2s_5_6(taps_imag_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_1_acc_nl[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl = (~ nor_491_tmp)
      & and_dcpl_209;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl = nor_491_tmp
      & and_dcpl_209;
  assign and_1537_nl = (((MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ MAC_2_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)) |
      MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp) & and_dcpl_976
      & and_dcpl_222;
  assign and_1541_nl = ((~ (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_2_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp) & (~((fsm_output[2])
      | MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp)) & and_dcpl_222;
  assign and_1544_nl = (((~ MAC_10_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp)
      & (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | MAC_10_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp) & and_dcpl_1054
      & and_dcpl_222;
  assign and_1548_nl = (MAC_10_ac_float_cctor_operator_1_ac_float_cctor_operator_1_nor_tmp
      | (~ (MAC_10_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & (~ MAC_10_ac_float_cctor_operator_ac_float_cctor_operator_nor_tmp) & and_dcpl_164
      & and_dcpl_222;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl = MUX_s_1_2_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_seb;
  assign and_2677_nl = (fsm_output[1]) & (~(((MAC_6_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_tmp[5])
      | (fsm_output[6])) & (fsm_output[0])));
  assign and_2678_nl = (fsm_output[1]) & (~((fsm_output[6]) & (fsm_output[0])));
  assign nor_751_nl = ~(and_dcpl_1363 | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_0
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_nand_5_itm));
  assign mux_567_nl = MUX_s_1_2_2(and_2677_nl, and_2678_nl, nor_751_nl);
  assign nor_807_nl = ~((fsm_output[6]) | (~ (fsm_output[0])));
  assign mux_568_nl = MUX_s_1_2_2(mux_567_nl, nor_807_nl, fsm_output[2]);
  assign nor_808_nl = ~((~((fsm_output[2:1]!=2'b10))) | (fsm_output[6]) | (fsm_output[0]));
  assign mux_569_nl = MUX_s_1_2_2(mux_568_nl, nor_808_nl, fsm_output[3]);
  assign nor_809_nl = ~((~ (fsm_output[1])) | (fsm_output[6]) | (fsm_output[0]));
  assign and_1285_nl = nor_98_cse & (~((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_218;
  assign and_1288_nl = nor_98_cse & (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_218;
  assign and_1291_nl = (~ (fsm_output[2])) & (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_218;
  assign and_1334_nl = nor_98_cse & (~((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      | MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_1450;
  assign and_1337_nl = nor_98_cse & (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_1450;
  assign and_1340_nl = (~ (fsm_output[2])) & (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_1450;
  assign and_942_nl = nor_98_cse & (~((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_1450;
  assign and_945_nl = nor_98_cse & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_1450;
  assign and_948_nl = (~ (fsm_output[2])) & (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_1450;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_1_nl
      = MUX1HOT_s_1_7_2((MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[4]), (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_4, (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[4]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0, {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_1_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_2_cse
      , and_1240_ssc , and_dcpl_574});
  assign and_1755_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_1_nl
      & (~ or_573_ssc) & (~ or_dcpl_577);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_4_nl
      = MUX1HOT_v_4_7_2((MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[3:0]), (MAC_2_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_19_3_0, (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_13_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[3:0]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1, {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_1_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_2_cse
      , and_1240_ssc , and_dcpl_574});
  assign nor_572_nl = ~(MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_4_nl,
      4'b1111, or_573_ssc));
  assign nor_571_nl = ~(MUX_v_4_2_2(nor_572_nl, 4'b1111, or_dcpl_577));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_2_nl
      = MUX1HOT_s_1_7_2((MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[4]), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_4, (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4]),
      (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[4]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0, {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_6_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_7_cse
      , and_1282_ssc , and_dcpl_624});
  assign and_1757_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_2_nl
      & (~ or_582_ssc) & (~ or_dcpl_578);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_5_nl
      = MUX1HOT_v_4_7_2((MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[3:0]), (MAC_3_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_17_3_0, (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[3:0]),
      (MAC_14_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_sdt[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[3:0]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1, {and_dcpl_189
      , and_dcpl_209 , and_dcpl_199 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_6_cse
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_and_7_cse
      , and_1282_ssc , and_dcpl_624});
  assign nor_570_nl = ~(MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_if_all_sign_1_mux1h_5_nl,
      4'b1111, or_582_ssc));
  assign nor_569_nl = ~(MUX_v_4_2_2(nor_570_nl, 4'b1111, or_dcpl_578));
  assign and_2681_nl = not_tmp_212 & (~ (fsm_output[6])) & (fsm_output[1]) & (~ (fsm_output[3]))
      & (fsm_output[0]) & (fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_2_nl
      = MUX_v_5_2_2((signext_5_4(~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_14_sva_6_0_rsp_2_rsp_1)),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_mux_1_cse, and_2681_nl);
  assign nl_z_out = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_2_nl)
      + 6'b000001;
  assign z_out = nl_z_out[5:0];
  assign and_2682_nl = not_tmp_212 & nor_501_cse & (fsm_output[2:0]==3'b111);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_3_nl
      = MUX_v_5_2_2((signext_5_4(~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0)),
      operator_i_e_1_lpi_1_dfm_mx0, and_2682_nl);
  assign nl_z_out_1 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_3_nl)
      + 6'b000001;
  assign z_out_1 = nl_z_out_1[5:0];
  assign and_2683_nl = nor_796_cse & (fsm_output[3:1]==3'b010);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_mux_1_nl
      = MUX_v_5_2_2((signext_5_4(~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[3:0]))),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1, and_2683_nl);
  assign nl_z_out_2 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_mux_1_nl)
      + 6'b000001;
  assign z_out_2 = nl_z_out_2[5:0];
  assign and_2684_nl = not_tmp_212 & (~((fsm_output[1:0]==2'b11))) & nor_501_cse
      & (fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl
      = MUX_v_5_2_2((signext_5_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_9_sva_rsp_1[3:0]))),
      ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_4 ,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_14_sva_3_0}),
      and_2684_nl);
  assign nl_z_out_3 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl)
      + 6'b000001;
  assign z_out_3 = nl_z_out_3[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_5_nl
      = MUX1HOT_s_1_4_2((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3])),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[5]),
      {and_1883_cse , and_1886_cse , and_1888_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_6_nl
      = MUX1HOT_s_1_4_2((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3])),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[5]),
      {and_1883_cse , and_1886_cse , and_1888_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_7_nl
      = MUX1HOT_v_5_4_2((signext_5_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[3:0]))),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_1_sva_6_0_rsp_2, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_10_itm_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_2_itm_rsp_1[4:0]),
      {and_1883_cse , and_1886_cse , and_1888_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_or_1_nl
      = (~((operator_ac_float_cctor_e_64_lpi_1_dfm[4]) | and_1883_cse)) | and_1888_cse
      | and_1893_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_8_nl
      = MUX1HOT_v_4_4_2(4'b0001, (~ (operator_ac_float_cctor_e_64_lpi_1_dfm[3:0])),
      (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0),
      (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0),
      {and_1883_cse , and_1886_cse , and_1888_cse , and_1893_cse});
  assign nl_acc_4_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_7_nl
      , (~ and_1883_cse)}) + conv_s2u_7_8({(~ and_1883_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_or_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux1h_8_nl
      , 1'b1});
  assign acc_4_nl = nl_acc_4_nl[7:0];
  assign z_out_4 = readslicef_8_7_1(acc_4_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_8_nl
      = MUX1HOT_s_1_4_2((~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2[3])),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0[5]),
      {and_1899_cse , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse
      , and_1886_cse , and_1888_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_9_nl
      = MUX1HOT_v_6_4_2((signext_6_4(~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_7_sva_6_0_rsp_2)),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_13_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_12_itm_5_0,
      {and_1899_cse , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse
      , and_1886_cse , and_1888_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_10_nl
      = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_4
      | and_1899_cse)) | and_1893_cse | and_1909_cse | and_1888_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_11_nl
      = and_1909_cse | and_1888_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_10_nl
      = MUX1HOT_v_4_4_2(4'b0001, (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0),
      (~ operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1), {and_1899_cse , and_1893_cse
      , and_1886_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_11_nl});
  assign nl_acc_5_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_9_nl
      , (~ and_1899_cse)}) + conv_s2u_7_8({(~ and_1899_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_10_nl
      , 1'b1});
  assign acc_5_nl = nl_acc_5_nl[7:0];
  assign z_out_5 = readslicef_8_7_1(acc_5_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_12_nl
      = and_dcpl_1780 | and_1909_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_13_nl
      = and_1925_cse | and_dcpl_1788;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_11_nl
      = MUX1HOT_v_6_3_2((signext_6_4(~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_8_sva_6_0_rsp_1[3:0]))),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_13_sva_rsp_1,
      {and_1899_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_13_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_14_nl
      = and_1909_cse | and_dcpl_1788;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_12_nl
      = MUX1HOT_v_4_4_2(4'b0001, (~ MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0),
      (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0), (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0),
      {and_1899_cse , and_dcpl_1780 , and_1925_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_or_14_nl});
  assign nl_acc_6_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_11_nl
      , (~ and_1899_cse)}) + conv_s2u_6_7({(~ and_1899_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux1h_12_nl
      , 1'b1});
  assign acc_6_nl = nl_acc_6_nl[6:0];
  assign z_out_6 = readslicef_7_6_1(acc_6_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_20_nl
      = MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0,
      {and_1883_cse , and_1888_cse , and_1886_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_21_nl
      = MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0[1]),
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_22_nl
      = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[4]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_0[0]),
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_23_nl
      = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_4_itm_5_0_rsp_1[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_15_itm_rsp_1_5_0_rsp_1,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_4_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[4])), (~ (operator_ac_float_cctor_e_14_lpi_1_dfm[4])),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_5_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_4_nl
      | and_1888_cse | and_1893_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_24_nl
      = MUX1HOT_v_4_4_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[3:0])), (~
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1),
      (~ (operator_ac_float_cctor_e_14_lpi_1_dfm[3:0])), (~ operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1),
      {and_1883_cse , and_1888_cse , and_1886_cse , and_1893_cse});
  assign nl_acc_7_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_20_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_22_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_23_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_24_nl
      , 1'b1});
  assign acc_7_nl = nl_acc_7_nl[7:0];
  assign z_out_7 = readslicef_8_7_1(acc_7_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_25_nl
      = MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_0,
      {and_1883_cse , and_1888_cse , and_1886_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl
      = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[5]),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_6_itm_5_0_rsp_1,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_13_sva_rsp_1_rsp_1[4:0]),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[4])), (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva[4])),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_6_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl
      | and_1888_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_26_nl
      = MUX1HOT_v_4_3_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[3:0])), (~
      operator_ac_float_cctor_m_61_lpi_1_dfm_rsp_1), (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_10_sva[3:0])),
      {and_1883_cse , and_1888_cse , and_1886_cse});
  assign nl_acc_8_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_25_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_26_nl
      , 1'b1});
  assign acc_8_nl = nl_acc_8_nl[7:0];
  assign z_out_8 = readslicef_8_7_1(acc_8_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl = MUX1HOT_s_1_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[5]),
      {and_1888_cse , and_1886_cse , and_1883_cse , and_1893_cse});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl = MUX1HOT_v_2_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[5:4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[5:4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[5:4]),
      {and_1888_cse , and_1886_cse , and_1883_cse , and_1893_cse});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl = MUX1HOT_v_4_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_2_itm_5_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]),
      {and_1888_cse , and_1886_cse , and_1883_cse , and_1893_cse});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_1_nl = MUX_s_1_2_2((~
      (operator_ac_float_cctor_e_3_lpi_1_dfm[4])), (~ (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[4])),
      and_1883_cse);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_nl
      = i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_1_nl | and_1888_cse
      | and_1893_cse;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl = MUX1HOT_v_4_4_2((~
      MAC_6_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0), (~ (operator_ac_float_cctor_e_3_lpi_1_dfm[3:0])),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[3:0])), (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0),
      {and_1888_cse , and_1886_cse , and_1883_cse , and_1893_cse});
  assign nl_acc_9_nl = ({i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl , 1'b1});
  assign acc_9_nl = nl_acc_9_nl[7:0];
  assign z_out_9 = readslicef_8_7_1(acc_9_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_27_nl
      = MUX1HOT_s_1_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0,
      {and_1883_cse , and_1888_cse , and_1886_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl
      = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0[1]),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_8_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[4]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0[0]),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_9_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_8_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1,
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[4])), (~ (operator_ac_float_cctor_e_29_lpi_1_dfm[4])),
      and_1886_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_7_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_6_nl
      | and_1888_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_28_nl
      = MUX1HOT_v_4_3_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[3:0])), (~
      operator_ac_float_cctor_m_62_lpi_1_dfm_rsp_1), (~ (operator_ac_float_cctor_e_29_lpi_1_dfm[3:0])),
      {and_1883_cse , and_1888_cse , and_1886_cse});
  assign nl_acc_10_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_27_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_9_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_28_nl
      , 1'b1});
  assign acc_10_nl = nl_acc_10_nl[7:0];
  assign z_out_10 = readslicef_8_7_1(acc_10_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_12_nl = and_dcpl_1857
      | and_dcpl_1860;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_0,
      {and_1925_cse , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_12_nl});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[5]),
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl
      = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_2_itm_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_14_sva_rsp_1[4:0]),
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl
      = (~((MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[4]) | and_dcpl_1860)) | and_1925_cse
      | and_1893_cse | and_1909_cse;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl = MUX1HOT_v_4_5_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_and_14_itm_3_0),
      (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_6_sva_1,
      (~ operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2), {and_1925_cse , and_1893_cse
      , and_dcpl_1857 , and_dcpl_1860 , and_1909_cse});
  assign nl_acc_11_nl = ({i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl
      , (~ and_dcpl_1860)}) + conv_s2u_7_8({(~ and_dcpl_1860) , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl , 1'b1});
  assign acc_11_nl = nl_acc_11_nl[7:0];
  assign z_out_11 = readslicef_8_7_1(acc_11_nl);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_13_nl = and_dcpl_1872
      | and_dcpl_1875;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[5]),
      {and_1925_cse , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_13_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse});
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[5]),
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl
      = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_4_itm_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_10_sva_rsp_1[4:0]),
      i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_cse);
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl
      = (~((MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[4]) | and_dcpl_1875)) | and_1925_cse
      | and_1909_cse | and_1893_cse;
  assign i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl = MUX1HOT_v_4_5_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_7_sva_1,
      (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_2_acc_itm_3_0), (~ operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2),
      {and_1925_cse , and_dcpl_1872 , and_dcpl_1875 , and_1909_cse , and_1893_cse});
  assign nl_acc_12_nl = ({i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl
      , (~ and_dcpl_1875)}) + conv_s2u_7_8({(~ and_dcpl_1875) , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl
      , i_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl , 1'b1});
  assign acc_12_nl = nl_acc_12_nl[7:0];
  assign z_out_12 = readslicef_8_7_1(acc_12_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_5_nl
      = MUX1HOT_s_1_4_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_0,
      {and_1886_cse , and_1893_cse , and_1888_cse , and_1883_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_6_nl
      = MUX1HOT_v_2_4_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[5:4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[5:4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_1,
      {and_1886_cse , and_1893_cse , and_1888_cse , and_1883_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_7_nl
      = MUX1HOT_v_4_4_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_14_itm_5_0[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_14_sva_6_0_rsp_2,
      {and_1886_cse , and_1893_cse , and_1888_cse , and_1883_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_22_nl
      = MUX_s_1_2_2((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[4])),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[4])), and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_or_1_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_22_nl
      | and_1893_cse | and_1888_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_8_nl
      = MUX1HOT_v_4_4_2((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_11_sva[3:0])),
      (~ operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1), (~ operator_ac_float_cctor_m_44_lpi_1_dfm_rsp_2),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[3:0])), {and_1886_cse , and_1893_cse
      , and_1888_cse , and_1883_cse});
  assign nl_acc_14_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_7_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_or_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_8_nl
      , 1'b1});
  assign acc_14_nl = nl_acc_14_nl[7:0];
  assign z_out_14 = readslicef_8_7_1(acc_14_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_4_nl
      = MUX1HOT_s_1_4_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1[5]),
      {and_1886_cse , and_1883_cse , and_1888_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_5_nl
      = MUX1HOT_v_6_4_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_11_sva_rsp_1_rsp_1,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1,
      {and_1886_cse , and_1883_cse , and_1888_cse , and_1893_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_23_nl
      = MUX_s_1_2_2((~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_4), (~
      (MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[4])), and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_1_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_23_nl
      | and_1888_cse | and_1893_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_3_nl
      = and_1888_cse | and_1893_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_6_nl
      = MUX1HOT_v_4_3_2((~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_3_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[3:0])), (~ MAC_5_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_3_acc_itm_3_0),
      {and_1886_cse , and_1883_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_3_nl});
  assign nl_acc_15_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_5_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_or_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux1h_6_nl
      , 1'b1});
  assign acc_15_nl = nl_acc_15_nl[7:0];
  assign z_out_15 = readslicef_8_7_1(acc_15_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl = and_dcpl_1939
      | and_dcpl_1942;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_14_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_0,
      {and_1893_cse , and_1925_cse , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[5]),
      and_1925_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl
      = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_4_itm_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_12_itm_rsp_1[4:0]),
      and_1925_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl
      = (~((MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[4]) | and_dcpl_1942)) | and_1893_cse
      | and_1925_cse;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl = MUX1HOT_v_4_4_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0),
      (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_6_sva_1,
      {and_1893_cse , and_1925_cse , and_dcpl_1939 , and_dcpl_1942});
  assign nl_acc_16_nl = ({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_14_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl
      , (~ and_dcpl_1942)}) + conv_s2u_7_8({(~ and_dcpl_1942) , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_6_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_15_nl , 1'b1});
  assign acc_16_nl = nl_acc_16_nl[7:0];
  assign z_out_16 = readslicef_8_7_1(acc_16_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_10_nl
      = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1[5]),
      and_1925_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_8_nl
      = (~((MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[4]) | and_dcpl_1962)) | and_1925_cse;
  assign and_2685_nl = and_dcpl_1740 & and_dcpl_1752 & (~((fsm_output[2]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_actual_max_shift_left_acc_psp_8_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_15_nl
      = MUX1HOT_v_4_3_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_8_sva_1,
      (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_12_sva_3_0),
      {and_2685_nl , and_dcpl_1962 , and_1925_cse});
  assign nl_acc_18_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_6_itm_rsp_1
      , (~ and_dcpl_1962)}) + conv_s2u_7_8({(~ and_dcpl_1962) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_15_nl
      , 1'b1});
  assign acc_18_nl = nl_acc_18_nl[7:0];
  assign z_out_18 = readslicef_8_7_1(acc_18_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_24_nl
      = MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0,
      (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2[3])),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_25_nl
      = MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1,
      (~ (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2[3])),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_26_nl
      = MUX_v_5_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2,
      (signext_5_4(~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_9_sva_6_0_rsp_2)),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_27_nl
      = MUX_v_5_2_2((~ operator_ac_float_cctor_e_65_lpi_1_dfm), 5'b00001, and_1883_cse);
  assign nl_acc_19_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_24_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_25_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_26_nl
      , (~ and_1883_cse)}) + conv_s2u_7_8({(~ and_1883_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_27_nl
      , 1'b1});
  assign acc_19_nl = nl_acc_19_nl[7:0];
  assign z_out_19 = readslicef_8_7_1(acc_19_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_0,
      and_2125_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl
      = ~((MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[4]) & and_2125_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl = MUX_v_4_2_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_5_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[3:0])), and_2125_cse);
  assign nl_acc_20_nl = ({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_8_itm_rsp_1
      , 1'b1}) + conv_s2u_7_8({1'b1 , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl , 1'b1});
  assign acc_20_nl = nl_acc_20_nl[7:0];
  assign z_out_20 = readslicef_8_7_1(acc_20_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_9_nl = and_dcpl_1995
      | and_dcpl_1998;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5]),
      {and_1893_cse , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_9_nl
      , and_1925_cse});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[5]),
      and_1925_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl
      = MUX_v_5_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_6_itm_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_14_itm_rsp_1[4:0]),
      and_1925_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl
      = (~((MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[4]) | and_dcpl_1998)) | and_1893_cse
      | and_1925_cse;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl = MUX1HOT_v_4_4_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_6_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_if_1_shift_r_7_sva_1,
      (~ operator_ac_float_cctor_m_50_lpi_1_dfm_rsp_1), {and_1893_cse , and_dcpl_1995
      , and_dcpl_1998 , and_1925_cse});
  assign nl_acc_21_nl = ({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_16_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_6_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl
      , (~ and_dcpl_1998)}) + conv_s2u_7_8({(~ and_dcpl_1998) , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_7_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_17_nl , 1'b1});
  assign acc_21_nl = nl_acc_21_nl[7:0];
  assign z_out_21 = readslicef_8_7_1(acc_21_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_28_nl
      = MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0,
      (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3])), and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_29_nl
      = MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1,
      (~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3])), and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_30_nl
      = MUX_v_5_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2,
      (signext_5_4(~ (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[3:0]))),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_0
      | and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_31_nl
      = MUX_v_4_2_2((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_12_sva_rsp_1),
      4'b0001, and_1883_cse);
  assign nl_acc_22_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_28_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_29_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_30_nl
      , (~ and_1883_cse)}) + conv_s2u_7_8({(~ and_1883_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_31_nl
      , 1'b1});
  assign acc_22_nl = nl_acc_22_nl[7:0];
  assign z_out_22 = readslicef_8_7_1(acc_22_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_32_nl
      = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_0,
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_33_nl
      = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1[1]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_1,
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_34_nl
      = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_1[0]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[4]),
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_35_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_1_sva_rsp_1_rsp_2,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_9_sva_6_0_rsp_2[3:0]),
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_36_nl
      = MUX_s_1_2_2((~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg[4])), and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_37_nl
      = MUX_v_4_2_2((~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_sva_4_0_rsp_1),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg[3:0])), and_2125_cse);
  assign nl_acc_23_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_32_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_33_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_34_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_35_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_36_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_37_nl
      , 1'b1});
  assign acc_23_nl = nl_acc_23_nl[7:0];
  assign z_out_23 = readslicef_8_7_1(acc_23_nl);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl = MUX1HOT_s_1_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_6,
      {and_1893_cse , and_1888_cse , and_1883_cse , and_1886_cse});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0[1]),
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl = MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[4]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_0[0]),
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl = MUX1HOT_v_4_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_mux1h_8_itm_rsp_1[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_itm_5_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_16_itm_rsp_1_5_0_rsp_1,
      {r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_5_cse_1 , and_1888_cse
      , and_1886_cse});
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl = MUX_s_1_2_2((~
      (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[4])), (~ (operator_ac_float_cctor_e_19_lpi_1_dfm[4])),
      and_1886_cse);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl
      = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux_7_nl | and_1893_cse
      | and_1888_cse;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl = MUX1HOT_v_4_4_2((~
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_7_sva_3_0),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_ls_4_0_13_sva_3_0),
      (~ (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[3:0])), (~ (operator_ac_float_cctor_e_19_lpi_1_dfm[3:0])),
      {and_1893_cse , and_1888_cse , and_1883_cse , and_1886_cse});
  assign nl_acc_25_nl = ({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_18_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_19_nl , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_20_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_21_nl , 1'b1})
      + conv_s2u_7_8({1'b1 , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_or_8_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_mux1h_22_nl , 1'b1});
  assign acc_25_nl = nl_acc_25_nl[7:0];
  assign z_out_25 = readslicef_8_7_1(acc_25_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_38_nl
      = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_0,
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3])),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_39_nl
      = MUX_v_6_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1,
      (signext_6_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_12_sva_rsp_1[3:0]))),
      and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl
      = ~(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_0 | and_1883_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_40_nl
      = MUX_v_4_2_2((~ operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_15_sva_4_0_rsp_1),
      4'b0001, and_1883_cse);
  assign nl_acc_26_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_38_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_39_nl
      , (~ and_1883_cse)}) + conv_s2u_7_8({(~ and_1883_cse) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_else_1_qelse_mux_40_nl
      , 1'b1});
  assign acc_26_nl = nl_acc_26_nl[7:0];
  assign z_out_26 = readslicef_8_7_1(acc_26_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_25_nl
      = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_6,
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_26_nl
      = MUX_v_2_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[5:4]),
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_27_nl
      = MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_itm_5_0[3:0]),
      and_2125_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_28_nl
      = MUX_v_5_2_2((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva),
      (~ MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg), and_2125_cse);
  assign nl_acc_27_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_25_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_26_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_27_nl
      , 1'b1}) + conv_s2u_7_8({1'b1 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_28_nl
      , 1'b1});
  assign acc_27_nl = nl_acc_27_nl[7:0];
  assign z_out_27 = readslicef_8_7_1(acc_27_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_3_nl
      = MUX_v_5_2_2((signext_5_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_acc_psp_11_sva_rsp_1[3:0]))),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2, and_2241_cse);
  assign nl_z_out_28 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_if_1_shift_r_mux_3_nl)
      + 6'b000001;
  assign z_out_28 = nl_z_out_28[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_4_nl
      = MUX_v_5_2_2((signext_5_4(~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_2_sva_rsp_1_rsp_1_rsp_1)),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_2_itm_5_0_rsp_1,
      and_2241_cse);
  assign nl_z_out_29 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_4_nl)
      + 6'b000001;
  assign z_out_29 = nl_z_out_29[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_5_nl
      = MUX_v_5_2_2((signext_5_4(~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_3_sva_rsp_1_rsp_2)),
      ({operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_4 , operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_6_0_rsp_1_3_0}),
      and_2241_cse);
  assign nl_z_out_30 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_if_1_shift_r_mux_5_nl)
      + 6'b000001;
  assign z_out_30 = nl_z_out_30[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_29_nl
      = MUX1HOT_v_5_4_2(({{4{ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6}},
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_6}),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_11_7, (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_10_6),
      (~ operator_ac_float_cctor_m_34_lpi_1_dfm_10_6), {and_1899_cse , and_1909_cse
      , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_30_nl
      = MUX1HOT_v_2_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[5:4]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_0, (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_5_4),
      (~ operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_0), {and_1899_cse , and_1909_cse
      , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_31_nl
      = MUX1HOT_v_4_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_mux1h_10_itm_5_0[3:0]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_12_sva_6_0_rsp_1[4:1]), (~
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_sva_3_0),
      (~ operator_ac_float_cctor_m_34_lpi_1_dfm_5_0_rsp_1), {and_1899_cse , and_1909_cse
      , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_2_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_8_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_2_nl,
      5'b11111, and_1899_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_9_nl
      = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0[1])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1)
      | and_1899_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[4])), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_0[0]),
      and_1909_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_1_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux_7_nl
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_1_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_32_nl
      = MUX1HOT_v_4_3_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_3_sva_rsp_1_rsp_1,
      4'b0001, {and_1899_cse , and_1909_cse , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_1_cse});
  assign nl_acc_31_nl = conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_29_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_30_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_31_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_cse})
      + conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_and_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_mux1h_32_nl
      , 1'b1});
  assign acc_31_nl = nl_acc_31_nl[12:0];
  assign z_out_33 = readslicef_13_12_1(acc_31_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_16_nl
      = MUX1HOT_v_5_3_2(({{4{ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0}},
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_0}),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_10_6),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_10_6),
      {and_1883_cse , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_17_nl
      = MUX1HOT_s_1_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_1,
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4[1])),
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4[1])),
      {and_1883_cse , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_18_nl
      = MUX1HOT_s_1_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[4]),
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_5_4[0])),
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_5_4[0])),
      {and_1883_cse , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_19_nl
      = MUX1HOT_v_4_3_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_8_sva_6_0_rsp_2[3:0]),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_sva_3_0),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_3_0),
      {and_1883_cse , and_2261_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_1_nl
      = MUX_v_5_2_2((~ MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg), 5'b00001, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_1_cse);
  assign nl_acc_32_nl = conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_16_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_17_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_19_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1})
      + conv_s2u_7_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_nor_1_cse_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_1_nl
      , 1'b1});
  assign acc_32_nl = nl_acc_32_nl[12:0];
  assign z_out_34 = readslicef_13_12_1(acc_32_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_20_nl
      = MUX1HOT_v_5_4_2(({{4{ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0}},
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_0}),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_11_7, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[11:7]),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_10_6),
      {and_1899_cse , and_1909_cse , and_2264_cse , and_2261_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_21_nl
      = MUX1HOT_s_1_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[5]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_0, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[6]),
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4[1])),
      {and_1899_cse , and_1909_cse , and_2264_cse , and_2261_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_22_nl
      = MUX1HOT_s_1_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[4]),
      operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_1, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[5]),
      (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_5_4[0])),
      {and_1899_cse , and_1909_cse , and_2264_cse , and_2261_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_23_nl
      = MUX1HOT_v_4_4_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_10_itm_rsp_1[3:0]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_11_sva_6_0_rsp_2[4:1]), (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_7_sva_mx0w1[4:1]),
      (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_sva_3_0),
      {and_1899_cse , and_1909_cse , and_2264_cse , and_2261_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_11_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_10_6,
      and_2264_cse);
  assign not_2701_nl = ~ and_2261_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_3_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_11_nl,
      not_2701_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_9_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_3_nl,
      5'b11111, and_1899_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_12_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0[1]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4[1]),
      and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_nor_3_nl
      = ~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_12_nl
      | and_1899_cse)) | and_2261_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_24_nl
      = MUX1HOT_s_1_3_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[4])), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_0[0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_5_4[0]),
      {and_1899_cse , and_1909_cse , and_2264_cse});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_4_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_24_nl
      & (~ and_2261_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_25_nl
      = MUX1HOT_v_4_4_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_2_sva_rsp_1_rsp_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_1_sva_3_0,
      4'b0001, {and_1899_cse , and_1909_cse , and_2264_cse , and_2261_cse});
  assign nl_acc_33_nl = conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_20_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_22_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_23_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_else_1_qelse_or_cse})
      + conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_and_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux1h_25_nl
      , 1'b1});
  assign acc_33_nl = nl_acc_33_nl[12:0];
  assign z_out_35 = readslicef_13_12_1(acc_33_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_13_nl
      = MUX_v_11_2_2((signext_11_7({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_12_itm_rsp_1})),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_8_sva_mx0w2[11:1]), and_2264_cse);
  assign not_2703_nl = ~ and_2264_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_10_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_10_6,
      5'b11111, not_2703_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4[1])
      | (~ and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_14_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[4])), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_5_4[0]),
      and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_15_nl
      = MUX_v_4_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_op2_21_11_3_sva_3_0,
      and_2264_cse);
  assign nl_acc_34_nl = conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_13_nl
      , (~ and_2264_cse)}) + conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_15_nl
      , 1'b1});
  assign acc_34_nl = nl_acc_34_nl[12:0];
  assign z_out_36 = readslicef_13_12_1(acc_34_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_16_nl
      = MUX_v_11_2_2((signext_11_7({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_mux1h_14_itm_rsp_1})),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_mx0w2[11:1]), and_2264_cse);
  assign not_2705_nl = ~ and_2264_cse;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_12_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_0,
      5'b11111, not_2705_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0[1])
      | (~ and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_17_nl
      = MUX_s_1_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[4])), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_0[0]),
      and_2264_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_18_nl
      = MUX_v_4_2_2((~ (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[3:0])), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_op2_21_11_5_sva_rsp_1_rsp_1,
      and_2264_cse);
  assign nl_acc_35_nl = conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_16_nl
      , (~ and_2264_cse)}) + conv_s2u_12_13({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_or_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_17_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_else_1_qelse_mux_18_nl
      , 1'b1});
  assign acc_35_nl = nl_acc_35_nl[12:0];
  assign z_out_37 = readslicef_13_12_1(acc_35_nl);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_7_nl =
      MUX_v_5_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_11_7, (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[11:7]),
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_8_nl =
      MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_0,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[6]), and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_9_nl =
      MUX_s_1_2_2(operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_1,
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[5]), and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_10_nl
      = MUX_v_4_2_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_10_sva_6_0_rsp_2[4:1]),
      (operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_5_sva_mx0w1[4:1]), and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_11_nl
      = MUX_v_5_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_0,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_10_6,
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_12_nl
      = MUX_v_2_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1[5:4]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_5_4,
      and_2317_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_13_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_1_op2_21_11_15_sva_rsp_1[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_sva_3_0,
      and_2317_cse);
  assign nl_z_out_38 = conv_s2u_11_12({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_7_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_8_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_9_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_10_nl})
      + conv_s2u_11_12({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_11_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_12_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_mux_13_nl});
  assign z_out_38 = nl_z_out_38[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_15_nl =
      MUX_v_12_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_9_sva[12:1]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_13_sva[12:1]),
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_16_nl =
      MUX_v_5_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_11_7,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6[5:1]),
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_17_nl =
      MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_0,
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_11_6[0]),
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_18_nl =
      MUX_v_2_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[5:4]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_5_4,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_19_nl =
      MUX_v_4_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_4_sva_6_0_rsp_1[3:0]),
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_22_itm_3_0,
      and_2326_cse);
  assign nl_z_out_39 = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_15_nl
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_16_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_17_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_18_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_19_nl});
  assign z_out_39 = nl_z_out_39[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_20_nl =
      MUX_v_12_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_3_sva[12:1]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_12_sva[12:1]),
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_21_nl =
      MUX_v_5_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_11_7,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_0,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_22_nl =
      MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_6,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_23_nl =
      MUX_v_2_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_5_4,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_24_nl =
      MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_add_r_12_1_6_sva_6_0_rsp_1_rsp_1,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_13_itm_rsp_1_3_0,
      and_2326_cse);
  assign nl_z_out_40 = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_20_nl
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_21_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_22_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_23_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_24_nl});
  assign z_out_40 = nl_z_out_40[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_25_nl =
      MUX_v_12_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_7_sva[12:1]),
      (ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_11_sva[12:1]),
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_26_nl =
      MUX_v_5_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_0,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_27_nl =
      MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_6,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_0,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_28_nl =
      MUX_v_2_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_5_4,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_0,
      and_2326_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_29_nl =
      MUX_v_4_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_10_itm_rsp_1_3_0,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_18_itm_rsp_1_rsp_1_rsp_1,
      and_2326_cse);
  assign nl_z_out_41 = ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_25_nl
      + ({ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_26_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_27_nl , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_28_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_mux_29_nl});
  assign z_out_41 = nl_z_out_41[11:0];
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_38_tmp
      = MUX_s_1_2_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[5]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[5]),
      and_2241_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_nl
      = ~(and_2241_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_38_tmp);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_3_nl =
      and_2241_cse & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_38_tmp);
  assign z_out_31 = MUX1HOT_v_5_3_2((operator_13_2_true_AC_TRN_AC_WRAP_1_rshift_psp_9_sva_6_0_rsp_1[4:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_itm_5_0[4:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_3_ls_4_0_sva, {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_3_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_38_tmp});
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc
      = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[1]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[5]),
      and_2241_cse);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_39_nl
      = MUX_s_1_2_2((ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_5_4[0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[4]),
      and_2241_cse);
  assign z_out_32_4 = MUX_s_1_2_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_39_nl,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva[4]), ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_1_nl
      = ~(and_2241_cse | ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc);
  assign ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_1_nl =
      and_2241_cse & (~ ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc);
  assign z_out_32_3_0 = MUX1HOT_v_4_3_2(ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_e_dif_acc_psp_11_sva_3_0,
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_2_acc_psp_14_sva_rsp_1[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ls_4_0_10_sva[3:0]),
      {ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_nor_1_nl
      , ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_and_1_nl ,
      ac_float_cctor_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_1_qelse_mux_41_ssc});

  function automatic  MUX1HOT_s_1_18_2;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [17:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    MUX1HOT_s_1_18_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_19_2;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [18:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    MUX1HOT_s_1_19_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_23_2;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [22:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    MUX1HOT_s_1_23_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_6_2;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [5:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    MUX1HOT_s_1_6_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_7_2;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [6:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_8_2;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [7:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    MUX1HOT_s_1_8_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_10_2;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [9:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    MUX1HOT_v_2_10_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_11_2;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [10:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    MUX1HOT_v_2_11_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_22_2;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [21:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    MUX1HOT_v_2_22_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_24_2;
    input [1:0] input_23;
    input [1:0] input_22;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [23:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    result = result | (input_22 & {2{sel[22]}});
    result = result | (input_23 & {2{sel[23]}});
    MUX1HOT_v_2_24_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_3_2;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [2:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    MUX1HOT_v_2_3_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_4_2;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [3:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    MUX1HOT_v_2_4_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_5_2;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [4:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    MUX1HOT_v_2_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_6_2;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [5:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    MUX1HOT_v_2_6_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_7_2;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [6:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    MUX1HOT_v_2_7_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_8_2;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [7:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    MUX1HOT_v_2_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_9_2;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [8:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    MUX1HOT_v_2_9_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_10_2;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [9:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    MUX1HOT_v_4_10_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_11_2;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [10:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    MUX1HOT_v_4_11_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_19_2;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [18:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    MUX1HOT_v_4_19_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_22_2;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [21:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    MUX1HOT_v_4_22_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_23_2;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [22:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    MUX1HOT_v_4_23_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_24_2;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [23:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    MUX1HOT_v_4_24_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_40_2;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [39:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    MUX1HOT_v_4_40_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_42_2;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [41:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    MUX1HOT_v_4_42_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_6_2;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [5:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    MUX1HOT_v_4_6_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_7_2;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [6:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    MUX1HOT_v_4_7_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_8_2;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [7:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    MUX1HOT_v_4_8_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_9_2;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [8:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    MUX1HOT_v_4_9_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_10_2;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [9:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    MUX1HOT_v_5_10_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_15_2;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [14:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    result = result | (input_13 & {5{sel[13]}});
    result = result | (input_14 & {5{sel[14]}});
    MUX1HOT_v_5_15_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_22_2;
    input [4:0] input_21;
    input [4:0] input_20;
    input [4:0] input_19;
    input [4:0] input_18;
    input [4:0] input_17;
    input [4:0] input_16;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [21:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    result = result | (input_13 & {5{sel[13]}});
    result = result | (input_14 & {5{sel[14]}});
    result = result | (input_15 & {5{sel[15]}});
    result = result | (input_16 & {5{sel[16]}});
    result = result | (input_17 & {5{sel[17]}});
    result = result | (input_18 & {5{sel[18]}});
    result = result | (input_19 & {5{sel[19]}});
    result = result | (input_20 & {5{sel[20]}});
    result = result | (input_21 & {5{sel[21]}});
    MUX1HOT_v_5_22_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_24_2;
    input [4:0] input_23;
    input [4:0] input_22;
    input [4:0] input_21;
    input [4:0] input_20;
    input [4:0] input_19;
    input [4:0] input_18;
    input [4:0] input_17;
    input [4:0] input_16;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [23:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    result = result | (input_13 & {5{sel[13]}});
    result = result | (input_14 & {5{sel[14]}});
    result = result | (input_15 & {5{sel[15]}});
    result = result | (input_16 & {5{sel[16]}});
    result = result | (input_17 & {5{sel[17]}});
    result = result | (input_18 & {5{sel[18]}});
    result = result | (input_19 & {5{sel[19]}});
    result = result | (input_20 & {5{sel[20]}});
    result = result | (input_21 & {5{sel[21]}});
    result = result | (input_22 & {5{sel[22]}});
    result = result | (input_23 & {5{sel[23]}});
    MUX1HOT_v_5_24_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_6_2;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [5:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    MUX1HOT_v_5_6_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_7_2;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [6:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    MUX1HOT_v_5_7_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_8_2;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [7:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    MUX1HOT_v_5_8_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_9_2;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [8:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    MUX1HOT_v_5_9_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_16_2;
    input [5:0] input_15;
    input [5:0] input_14;
    input [5:0] input_13;
    input [5:0] input_12;
    input [5:0] input_11;
    input [5:0] input_10;
    input [5:0] input_9;
    input [5:0] input_8;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [15:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    result = result | (input_8 & {6{sel[8]}});
    result = result | (input_9 & {6{sel[9]}});
    result = result | (input_10 & {6{sel[10]}});
    result = result | (input_11 & {6{sel[11]}});
    result = result | (input_12 & {6{sel[12]}});
    result = result | (input_13 & {6{sel[13]}});
    result = result | (input_14 & {6{sel[14]}});
    result = result | (input_15 & {6{sel[15]}});
    MUX1HOT_v_6_16_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_3_2;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [2:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    MUX1HOT_v_6_3_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_4_2;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [3:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    MUX1HOT_v_6_4_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_5_2;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [4:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    MUX1HOT_v_6_5_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_6_2;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [5:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    MUX1HOT_v_6_6_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_7_2;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [6:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    MUX1HOT_v_6_7_2 = result;
  end
  endfunction


  function automatic [5:0] MUX1HOT_v_6_8_2;
    input [5:0] input_7;
    input [5:0] input_6;
    input [5:0] input_5;
    input [5:0] input_4;
    input [5:0] input_3;
    input [5:0] input_2;
    input [5:0] input_1;
    input [5:0] input_0;
    input [7:0] sel;
    reg [5:0] result;
  begin
    result = input_0 & {6{sel[0]}};
    result = result | (input_1 & {6{sel[1]}});
    result = result | (input_2 & {6{sel[2]}});
    result = result | (input_3 & {6{sel[3]}});
    result = result | (input_4 & {6{sel[4]}});
    result = result | (input_5 & {6{sel[5]}});
    result = result | (input_6 & {6{sel[6]}});
    result = result | (input_7 & {6{sel[7]}});
    MUX1HOT_v_6_8_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [11:0] MUX_v_12_2_2;
    input [11:0] input_0;
    input [11:0] input_1;
    input  sel;
    reg [11:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_12_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [11:0] readslicef_13_12_1;
    input [12:0] vector;
    reg [12:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_13_12_1 = tmp[11:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [5:0] readslicef_7_6_1;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_7_6_1 = tmp[5:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [10:0] signext_11_7;
    input [6:0] vector;
  begin
    signext_11_7= {{4{vector[6]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_4;
    input [3:0] vector;
  begin
    signext_5_4= {{1{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] signext_6_4;
    input [3:0] vector;
  begin
    signext_6_4= {{2{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [11:0] conv_s2s_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2s_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2u_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2u_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [7:0] conv_s2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_7_13 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_13 = {{6{vector[6]}}, vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [12:0] conv_s2u_12_13 ;
    input [11:0]  vector ;
  begin
    conv_s2u_12_13 = {vector[11], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_4_7 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_7 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_real_m_rsc_dat, input_real_m_triosy_lz, input_real_e_rsc_dat, input_real_e_triosy_lz,
      input_imag_m_rsc_dat, input_imag_m_triosy_lz, input_imag_e_rsc_dat, input_imag_e_triosy_lz,
      taps_real_m_rsc_dat, taps_real_m_triosy_lz, taps_real_e_rsc_dat, taps_real_e_triosy_lz,
      taps_imag_m_rsc_dat, taps_imag_m_triosy_lz, taps_imag_e_rsc_dat, taps_imag_e_triosy_lz,
      return_real_m_rsc_dat, return_real_m_triosy_lz, return_real_e_rsc_dat, return_real_e_triosy_lz,
      return_imag_m_rsc_dat, return_imag_m_triosy_lz, return_imag_e_rsc_dat, return_imag_e_triosy_lz
);
  input clk;
  input rst;
  input [10:0] input_real_m_rsc_dat;
  output input_real_m_triosy_lz;
  input [4:0] input_real_e_rsc_dat;
  output input_real_e_triosy_lz;
  input [10:0] input_imag_m_rsc_dat;
  output input_imag_m_triosy_lz;
  input [4:0] input_imag_e_rsc_dat;
  output input_imag_e_triosy_lz;
  input [175:0] taps_real_m_rsc_dat;
  output taps_real_m_triosy_lz;
  input [79:0] taps_real_e_rsc_dat;
  output taps_real_e_triosy_lz;
  input [175:0] taps_imag_m_rsc_dat;
  output taps_imag_m_triosy_lz;
  input [79:0] taps_imag_e_rsc_dat;
  output taps_imag_e_triosy_lz;
  output [10:0] return_real_m_rsc_dat;
  output return_real_m_triosy_lz;
  output [4:0] return_real_e_rsc_dat;
  output return_real_e_triosy_lz;
  output [10:0] return_imag_m_rsc_dat;
  output return_imag_m_triosy_lz;
  output [4:0] return_imag_e_rsc_dat;
  output return_imag_e_triosy_lz;


  // Interconnect Declarations
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;


  // Interconnect Declarations for Component Instantiations 
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_1 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_2 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_3 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_4 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_5 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_6 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_7 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_8 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_9 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_10 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_11 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_12 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_13 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_14 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_15 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_16 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_17 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_18 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_19 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_20 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_21 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_22 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_23 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_24 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_25 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_26 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_27 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_28 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_29 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_30 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_31 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_32 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_33 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_34 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_35 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_36 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_37 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_38 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_39 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_40 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_41 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_42 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_43 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_44 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_45 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_46 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_47 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_48 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_49 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_50 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_51 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_52 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_53 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_54 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_55 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_56 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_57 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_58 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_59 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_60 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_61 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_62 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_63 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn)
    );
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .input_real_m_rsc_dat(input_real_m_rsc_dat),
      .input_real_m_triosy_lz(input_real_m_triosy_lz),
      .input_real_e_rsc_dat(input_real_e_rsc_dat),
      .input_real_e_triosy_lz(input_real_e_triosy_lz),
      .input_imag_m_rsc_dat(input_imag_m_rsc_dat),
      .input_imag_m_triosy_lz(input_imag_m_triosy_lz),
      .input_imag_e_rsc_dat(input_imag_e_rsc_dat),
      .input_imag_e_triosy_lz(input_imag_e_triosy_lz),
      .taps_real_m_rsc_dat(taps_real_m_rsc_dat),
      .taps_real_m_triosy_lz(taps_real_m_triosy_lz),
      .taps_real_e_rsc_dat(taps_real_e_rsc_dat),
      .taps_real_e_triosy_lz(taps_real_e_triosy_lz),
      .taps_imag_m_rsc_dat(taps_imag_m_rsc_dat),
      .taps_imag_m_triosy_lz(taps_imag_m_triosy_lz),
      .taps_imag_e_rsc_dat(taps_imag_e_rsc_dat),
      .taps_imag_e_triosy_lz(taps_imag_e_triosy_lz),
      .return_real_m_rsc_dat(return_real_m_rsc_dat),
      .return_real_m_triosy_lz(return_real_m_triosy_lz),
      .return_real_e_rsc_dat(return_real_e_rsc_dat),
      .return_real_e_triosy_lz(return_real_e_triosy_lz),
      .return_imag_m_rsc_dat(return_imag_m_rsc_dat),
      .return_imag_m_triosy_lz(return_imag_m_triosy_lz),
      .return_imag_e_rsc_dat(return_imag_e_rsc_dat),
      .return_imag_e_triosy_lz(return_imag_e_triosy_lz),
      .MAC_1_leading_sign_18_1_1_0_cmp_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn)
    );
endmodule



