
//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/ccs_out_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_out_v1 (dat, idat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output   [width-1:0] dat;
  input    [width-1:0] idat;

  wire     [width-1:0] dat;

  assign dat = idat;

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_io_sync_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_io_sync_v2 (ld, lz);
    parameter valid = 0;

    input  ld;
    output lz;

    wire   lz;

    assign lz = ld;

endmodule


//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_r_beh_v5.v 
module mgc_shift_r_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_u(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_u(a,s,1'b0);
     end
   endgenerate

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/leading_sign_13_1_1_0_fbd6b6484e0226fdfa7c7e6838ce99f45fe9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:36 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_13_1_1_0
// ------------------------------------------------------------------


module leading_sign_13_1_1_0 (
  mantissa, all_same, rtn
);
  input [12:0] mantissa;
  output all_same;
  output [3:0] rtn;


  // Interconnect Declarations
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire [11:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0;
  wire c_h_1_2;
  wire c_h_1_4;

  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl;
  wire[1:0] r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl;
  wire r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl;

  // Interconnect Declarations for Component Instantiations 
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0 = (mantissa[11:0])
      ^ (signext_12_1(~ (mantissa[12])));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[9:8]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1 =
      (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11:10]==2'b11);
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7:6]==2'b11);
  assign c_h_1_2 = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[5:4]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3:2]==2'b11);
  assign c_h_1_4 = c_h_1_2 & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4
      = (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[1:0]==2'b11)
      & r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1 &
      c_h_1_4;
  assign all_same = r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      = (c_h_1_2 & (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_18_3_sdt_3))
      | r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4;
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl = ~(r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_1
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_26_2_sdt_1
      | (~ c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl = ~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[11])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[10:9]!=2'b10))
      & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[7])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[6:5]!=2'b10))))
      & c_h_1_2)) & (~((~((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[3])
      & ((r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_xor_11_0[2:1]!=2'b10))))
      & c_h_1_4)));
  assign r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl
      = ~(MUX_v_2_2_2(({r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nand_2_nl}), 2'b11,
      r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_wrs_c_32_4_sdt_4));
  assign rtn = {c_h_1_4 , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_or_1_nl
      , r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_r_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_all_sign_1_nor_nl};

  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [11:0] signext_12_1;
    input  vector;
  begin
    signext_12_1= {{11{vector}}, vector};
  end
  endfunction

endmodule




//------> /eda/mentor/Siemens_EDA/Catapult_Synthesis_2023.1_2/Mgc_home/pkgs/siflibs/mgc_shift_br_beh_v5.v 
module mgc_shift_br_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
     if (signd_a)
     begin: SGNED
       assign z = fshr_s(a,s,a[width_a-1]);
     end
     else
     begin: UNSGNED
       assign z = fshr_s(a,s,1'b0);
     end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift right - unsigned shift argument
   function [width_z-1:0] fshr_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = signd_a ? width_a : width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg signed [len-1:0] result;
      reg signed [len-1:0] result_t;
      begin
        result_t = $signed( {(len){sbit}} );
        result_t[width_a-1:0] = arg1;
        result = result_t >>> arg2;
        fshr_u =  result[olen-1:0];
      end
   endfunction // fshr_u

   //Shift right - signed shift argument
   function [width_z-1:0] fshr_s;
     input [width_a-1:0] arg1;
     input [width_s-1:0] arg2;
     input sbit;
     begin
       if ( arg2[width_s-1] == 1'b0 )
       begin
         fshr_s = fshr_u(arg1, arg2, sbit);
       end
       else
       begin
         fshr_s = fshl_u_1({arg1, 1'b0},~arg2, sbit);
       end
     end
   endfunction 

endmodule

//------> ../td_ccore_solutions/leading_sign_18_1_1_0_7b2153b3b691fe1ab68d43c72c494a7b6845_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Tue Apr 22 14:20:37 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    leading_sign_18_1_1_0
// ------------------------------------------------------------------


module leading_sign_18_1_1_0 (
  mantissa, all_same, rtn
);
  input [17:0] mantissa;
  output all_same;
  output [4:0] rtn;


  // Interconnect Declarations
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1;
  wire [16:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0;
  wire c_h_1_2;
  wire c_h_1_5;
  wire c_h_1_6;
  wire c_h_1_7;

  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl;

  // Interconnect Declarations for Component Instantiations 
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0
      = (mantissa[16:0]) ^ (signext_17_1(~ (mantissa[17])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[14:13]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16:15]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12:11]==2'b11);
  assign c_h_1_2 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[10:9]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[6:5]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8:7]==2'b11);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4:3]==2'b11);
  assign c_h_1_5 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[2:1]==2'b11)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      & c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[0])
      & c_h_1_7;
  assign all_same = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      = c_h_1_6 & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_42_4_sdt_4);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      = c_h_1_2 & (c_h_1_5 | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_18_3_sdt_3))
      & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_14_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_6_2_sdt_2))
      & (~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_1
      & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_34_2_sdt_1
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_26_2_sdt_2))))
      & c_h_1_6)) & (~ c_h_1_7);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl
      = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[16])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[15:14]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[12])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[11:10]!=2'b10))))
      & c_h_1_2)) & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[8])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[7:6]!=2'b10))
      & (~((~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[4])
      & ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_xor_16_0[3:2]!=2'b10))))
      & c_h_1_5)))) & c_h_1_6)) & (~ c_h_1_7)) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_wrs_c_48_5_sdt_5;
  assign rtn = {c_h_1_7 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_1_nl};

  function automatic [16:0] signext_17_1;
    input  vector;
  begin
    signext_17_1= {{16{vector}}, vector};
  end
  endfunction

endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2023.1_2/1049935 Production Release
//  HLS Date:       Sat Jun 10 10:53:51 PDT 2023
// 
//  Generated by:   ajh9498@hansolo.poly.edu
//  Generated date: Thu Apr 24 04:43:26 2025
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    fir_core_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module fir_core_core_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [8:0] fsm_output;
  reg [8:0] fsm_output;


  // FSM State Type Declaration for fir_core_core_fsm_1
  parameter
    main_C_0 = 9'd0,
    main_C_1 = 9'd1,
    main_C_2 = 9'd2,
    main_C_3 = 9'd3,
    main_C_4 = 9'd4,
    main_C_5 = 9'd5,
    main_C_6 = 9'd6,
    main_C_7 = 9'd7,
    main_C_8 = 9'd8,
    main_C_9 = 9'd9,
    main_C_10 = 9'd10,
    main_C_11 = 9'd11,
    main_C_12 = 9'd12,
    main_C_13 = 9'd13,
    main_C_14 = 9'd14,
    main_C_15 = 9'd15,
    main_C_16 = 9'd16,
    main_C_17 = 9'd17,
    main_C_18 = 9'd18,
    main_C_19 = 9'd19,
    main_C_20 = 9'd20,
    main_C_21 = 9'd21,
    main_C_22 = 9'd22,
    main_C_23 = 9'd23,
    main_C_24 = 9'd24,
    main_C_25 = 9'd25,
    main_C_26 = 9'd26,
    main_C_27 = 9'd27,
    main_C_28 = 9'd28,
    main_C_29 = 9'd29,
    main_C_30 = 9'd30,
    main_C_31 = 9'd31,
    main_C_32 = 9'd32,
    main_C_33 = 9'd33,
    main_C_34 = 9'd34,
    main_C_35 = 9'd35,
    main_C_36 = 9'd36,
    main_C_37 = 9'd37,
    main_C_38 = 9'd38,
    main_C_39 = 9'd39,
    main_C_40 = 9'd40,
    main_C_41 = 9'd41,
    main_C_42 = 9'd42,
    main_C_43 = 9'd43,
    main_C_44 = 9'd44,
    main_C_45 = 9'd45,
    main_C_46 = 9'd46,
    main_C_47 = 9'd47,
    main_C_48 = 9'd48,
    main_C_49 = 9'd49,
    main_C_50 = 9'd50,
    main_C_51 = 9'd51,
    main_C_52 = 9'd52,
    main_C_53 = 9'd53,
    main_C_54 = 9'd54,
    main_C_55 = 9'd55,
    main_C_56 = 9'd56,
    main_C_57 = 9'd57,
    main_C_58 = 9'd58,
    main_C_59 = 9'd59,
    main_C_60 = 9'd60,
    main_C_61 = 9'd61,
    main_C_62 = 9'd62,
    main_C_63 = 9'd63,
    main_C_64 = 9'd64,
    main_C_65 = 9'd65,
    main_C_66 = 9'd66,
    main_C_67 = 9'd67,
    main_C_68 = 9'd68,
    main_C_69 = 9'd69,
    main_C_70 = 9'd70,
    main_C_71 = 9'd71,
    main_C_72 = 9'd72,
    main_C_73 = 9'd73,
    main_C_74 = 9'd74,
    main_C_75 = 9'd75,
    main_C_76 = 9'd76,
    main_C_77 = 9'd77,
    main_C_78 = 9'd78,
    main_C_79 = 9'd79,
    main_C_80 = 9'd80,
    main_C_81 = 9'd81,
    main_C_82 = 9'd82,
    main_C_83 = 9'd83,
    main_C_84 = 9'd84,
    main_C_85 = 9'd85,
    main_C_86 = 9'd86,
    main_C_87 = 9'd87,
    main_C_88 = 9'd88,
    main_C_89 = 9'd89,
    main_C_90 = 9'd90,
    main_C_91 = 9'd91,
    main_C_92 = 9'd92,
    main_C_93 = 9'd93,
    main_C_94 = 9'd94,
    main_C_95 = 9'd95,
    main_C_96 = 9'd96,
    main_C_97 = 9'd97,
    main_C_98 = 9'd98,
    main_C_99 = 9'd99,
    main_C_100 = 9'd100,
    main_C_101 = 9'd101,
    main_C_102 = 9'd102,
    main_C_103 = 9'd103,
    main_C_104 = 9'd104,
    main_C_105 = 9'd105,
    main_C_106 = 9'd106,
    main_C_107 = 9'd107,
    main_C_108 = 9'd108,
    main_C_109 = 9'd109,
    main_C_110 = 9'd110,
    main_C_111 = 9'd111,
    main_C_112 = 9'd112,
    main_C_113 = 9'd113,
    main_C_114 = 9'd114,
    main_C_115 = 9'd115,
    main_C_116 = 9'd116,
    main_C_117 = 9'd117,
    main_C_118 = 9'd118,
    main_C_119 = 9'd119,
    main_C_120 = 9'd120,
    main_C_121 = 9'd121,
    main_C_122 = 9'd122,
    main_C_123 = 9'd123,
    main_C_124 = 9'd124,
    main_C_125 = 9'd125,
    main_C_126 = 9'd126,
    main_C_127 = 9'd127,
    main_C_128 = 9'd128,
    main_C_129 = 9'd129,
    main_C_130 = 9'd130,
    main_C_131 = 9'd131,
    main_C_132 = 9'd132,
    main_C_133 = 9'd133,
    main_C_134 = 9'd134,
    main_C_135 = 9'd135,
    main_C_136 = 9'd136,
    main_C_137 = 9'd137,
    main_C_138 = 9'd138,
    main_C_139 = 9'd139,
    main_C_140 = 9'd140,
    main_C_141 = 9'd141,
    main_C_142 = 9'd142,
    main_C_143 = 9'd143,
    main_C_144 = 9'd144,
    main_C_145 = 9'd145,
    main_C_146 = 9'd146,
    main_C_147 = 9'd147,
    main_C_148 = 9'd148,
    main_C_149 = 9'd149,
    main_C_150 = 9'd150,
    main_C_151 = 9'd151,
    main_C_152 = 9'd152,
    main_C_153 = 9'd153,
    main_C_154 = 9'd154,
    main_C_155 = 9'd155,
    main_C_156 = 9'd156,
    main_C_157 = 9'd157,
    main_C_158 = 9'd158,
    main_C_159 = 9'd159,
    main_C_160 = 9'd160,
    main_C_161 = 9'd161,
    main_C_162 = 9'd162,
    main_C_163 = 9'd163,
    main_C_164 = 9'd164,
    main_C_165 = 9'd165,
    main_C_166 = 9'd166,
    main_C_167 = 9'd167,
    main_C_168 = 9'd168,
    main_C_169 = 9'd169,
    main_C_170 = 9'd170,
    main_C_171 = 9'd171,
    main_C_172 = 9'd172,
    main_C_173 = 9'd173,
    main_C_174 = 9'd174,
    main_C_175 = 9'd175,
    main_C_176 = 9'd176,
    main_C_177 = 9'd177,
    main_C_178 = 9'd178,
    main_C_179 = 9'd179,
    main_C_180 = 9'd180,
    main_C_181 = 9'd181,
    main_C_182 = 9'd182,
    main_C_183 = 9'd183,
    main_C_184 = 9'd184,
    main_C_185 = 9'd185,
    main_C_186 = 9'd186,
    main_C_187 = 9'd187,
    main_C_188 = 9'd188,
    main_C_189 = 9'd189,
    main_C_190 = 9'd190,
    main_C_191 = 9'd191,
    main_C_192 = 9'd192,
    main_C_193 = 9'd193,
    main_C_194 = 9'd194,
    main_C_195 = 9'd195,
    main_C_196 = 9'd196,
    main_C_197 = 9'd197,
    main_C_198 = 9'd198,
    main_C_199 = 9'd199,
    main_C_200 = 9'd200,
    main_C_201 = 9'd201,
    main_C_202 = 9'd202,
    main_C_203 = 9'd203,
    main_C_204 = 9'd204,
    main_C_205 = 9'd205,
    main_C_206 = 9'd206,
    main_C_207 = 9'd207,
    main_C_208 = 9'd208,
    main_C_209 = 9'd209,
    main_C_210 = 9'd210,
    main_C_211 = 9'd211,
    main_C_212 = 9'd212,
    main_C_213 = 9'd213,
    main_C_214 = 9'd214,
    main_C_215 = 9'd215,
    main_C_216 = 9'd216,
    main_C_217 = 9'd217,
    main_C_218 = 9'd218,
    main_C_219 = 9'd219,
    main_C_220 = 9'd220,
    main_C_221 = 9'd221,
    main_C_222 = 9'd222,
    main_C_223 = 9'd223,
    main_C_224 = 9'd224,
    main_C_225 = 9'd225,
    main_C_226 = 9'd226,
    main_C_227 = 9'd227,
    main_C_228 = 9'd228,
    main_C_229 = 9'd229,
    main_C_230 = 9'd230,
    main_C_231 = 9'd231,
    main_C_232 = 9'd232,
    main_C_233 = 9'd233,
    main_C_234 = 9'd234,
    main_C_235 = 9'd235,
    main_C_236 = 9'd236,
    main_C_237 = 9'd237,
    main_C_238 = 9'd238,
    main_C_239 = 9'd239,
    main_C_240 = 9'd240,
    main_C_241 = 9'd241,
    main_C_242 = 9'd242,
    main_C_243 = 9'd243,
    main_C_244 = 9'd244,
    main_C_245 = 9'd245,
    main_C_246 = 9'd246,
    main_C_247 = 9'd247,
    main_C_248 = 9'd248,
    main_C_249 = 9'd249,
    main_C_250 = 9'd250,
    main_C_251 = 9'd251,
    main_C_252 = 9'd252,
    main_C_253 = 9'd253,
    main_C_254 = 9'd254,
    main_C_255 = 9'd255,
    main_C_256 = 9'd256,
    main_C_257 = 9'd257,
    main_C_258 = 9'd258;

  reg [8:0] state_var;
  reg [8:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : fir_core_core_fsm_1
    case (state_var)
      main_C_1 : begin
        fsm_output = 9'b000000001;
        state_var_NS = main_C_2;
      end
      main_C_2 : begin
        fsm_output = 9'b000000010;
        state_var_NS = main_C_3;
      end
      main_C_3 : begin
        fsm_output = 9'b000000011;
        state_var_NS = main_C_4;
      end
      main_C_4 : begin
        fsm_output = 9'b000000100;
        state_var_NS = main_C_5;
      end
      main_C_5 : begin
        fsm_output = 9'b000000101;
        state_var_NS = main_C_6;
      end
      main_C_6 : begin
        fsm_output = 9'b000000110;
        state_var_NS = main_C_7;
      end
      main_C_7 : begin
        fsm_output = 9'b000000111;
        state_var_NS = main_C_8;
      end
      main_C_8 : begin
        fsm_output = 9'b000001000;
        state_var_NS = main_C_9;
      end
      main_C_9 : begin
        fsm_output = 9'b000001001;
        state_var_NS = main_C_10;
      end
      main_C_10 : begin
        fsm_output = 9'b000001010;
        state_var_NS = main_C_11;
      end
      main_C_11 : begin
        fsm_output = 9'b000001011;
        state_var_NS = main_C_12;
      end
      main_C_12 : begin
        fsm_output = 9'b000001100;
        state_var_NS = main_C_13;
      end
      main_C_13 : begin
        fsm_output = 9'b000001101;
        state_var_NS = main_C_14;
      end
      main_C_14 : begin
        fsm_output = 9'b000001110;
        state_var_NS = main_C_15;
      end
      main_C_15 : begin
        fsm_output = 9'b000001111;
        state_var_NS = main_C_16;
      end
      main_C_16 : begin
        fsm_output = 9'b000010000;
        state_var_NS = main_C_17;
      end
      main_C_17 : begin
        fsm_output = 9'b000010001;
        state_var_NS = main_C_18;
      end
      main_C_18 : begin
        fsm_output = 9'b000010010;
        state_var_NS = main_C_19;
      end
      main_C_19 : begin
        fsm_output = 9'b000010011;
        state_var_NS = main_C_20;
      end
      main_C_20 : begin
        fsm_output = 9'b000010100;
        state_var_NS = main_C_21;
      end
      main_C_21 : begin
        fsm_output = 9'b000010101;
        state_var_NS = main_C_22;
      end
      main_C_22 : begin
        fsm_output = 9'b000010110;
        state_var_NS = main_C_23;
      end
      main_C_23 : begin
        fsm_output = 9'b000010111;
        state_var_NS = main_C_24;
      end
      main_C_24 : begin
        fsm_output = 9'b000011000;
        state_var_NS = main_C_25;
      end
      main_C_25 : begin
        fsm_output = 9'b000011001;
        state_var_NS = main_C_26;
      end
      main_C_26 : begin
        fsm_output = 9'b000011010;
        state_var_NS = main_C_27;
      end
      main_C_27 : begin
        fsm_output = 9'b000011011;
        state_var_NS = main_C_28;
      end
      main_C_28 : begin
        fsm_output = 9'b000011100;
        state_var_NS = main_C_29;
      end
      main_C_29 : begin
        fsm_output = 9'b000011101;
        state_var_NS = main_C_30;
      end
      main_C_30 : begin
        fsm_output = 9'b000011110;
        state_var_NS = main_C_31;
      end
      main_C_31 : begin
        fsm_output = 9'b000011111;
        state_var_NS = main_C_32;
      end
      main_C_32 : begin
        fsm_output = 9'b000100000;
        state_var_NS = main_C_33;
      end
      main_C_33 : begin
        fsm_output = 9'b000100001;
        state_var_NS = main_C_34;
      end
      main_C_34 : begin
        fsm_output = 9'b000100010;
        state_var_NS = main_C_35;
      end
      main_C_35 : begin
        fsm_output = 9'b000100011;
        state_var_NS = main_C_36;
      end
      main_C_36 : begin
        fsm_output = 9'b000100100;
        state_var_NS = main_C_37;
      end
      main_C_37 : begin
        fsm_output = 9'b000100101;
        state_var_NS = main_C_38;
      end
      main_C_38 : begin
        fsm_output = 9'b000100110;
        state_var_NS = main_C_39;
      end
      main_C_39 : begin
        fsm_output = 9'b000100111;
        state_var_NS = main_C_40;
      end
      main_C_40 : begin
        fsm_output = 9'b000101000;
        state_var_NS = main_C_41;
      end
      main_C_41 : begin
        fsm_output = 9'b000101001;
        state_var_NS = main_C_42;
      end
      main_C_42 : begin
        fsm_output = 9'b000101010;
        state_var_NS = main_C_43;
      end
      main_C_43 : begin
        fsm_output = 9'b000101011;
        state_var_NS = main_C_44;
      end
      main_C_44 : begin
        fsm_output = 9'b000101100;
        state_var_NS = main_C_45;
      end
      main_C_45 : begin
        fsm_output = 9'b000101101;
        state_var_NS = main_C_46;
      end
      main_C_46 : begin
        fsm_output = 9'b000101110;
        state_var_NS = main_C_47;
      end
      main_C_47 : begin
        fsm_output = 9'b000101111;
        state_var_NS = main_C_48;
      end
      main_C_48 : begin
        fsm_output = 9'b000110000;
        state_var_NS = main_C_49;
      end
      main_C_49 : begin
        fsm_output = 9'b000110001;
        state_var_NS = main_C_50;
      end
      main_C_50 : begin
        fsm_output = 9'b000110010;
        state_var_NS = main_C_51;
      end
      main_C_51 : begin
        fsm_output = 9'b000110011;
        state_var_NS = main_C_52;
      end
      main_C_52 : begin
        fsm_output = 9'b000110100;
        state_var_NS = main_C_53;
      end
      main_C_53 : begin
        fsm_output = 9'b000110101;
        state_var_NS = main_C_54;
      end
      main_C_54 : begin
        fsm_output = 9'b000110110;
        state_var_NS = main_C_55;
      end
      main_C_55 : begin
        fsm_output = 9'b000110111;
        state_var_NS = main_C_56;
      end
      main_C_56 : begin
        fsm_output = 9'b000111000;
        state_var_NS = main_C_57;
      end
      main_C_57 : begin
        fsm_output = 9'b000111001;
        state_var_NS = main_C_58;
      end
      main_C_58 : begin
        fsm_output = 9'b000111010;
        state_var_NS = main_C_59;
      end
      main_C_59 : begin
        fsm_output = 9'b000111011;
        state_var_NS = main_C_60;
      end
      main_C_60 : begin
        fsm_output = 9'b000111100;
        state_var_NS = main_C_61;
      end
      main_C_61 : begin
        fsm_output = 9'b000111101;
        state_var_NS = main_C_62;
      end
      main_C_62 : begin
        fsm_output = 9'b000111110;
        state_var_NS = main_C_63;
      end
      main_C_63 : begin
        fsm_output = 9'b000111111;
        state_var_NS = main_C_64;
      end
      main_C_64 : begin
        fsm_output = 9'b001000000;
        state_var_NS = main_C_65;
      end
      main_C_65 : begin
        fsm_output = 9'b001000001;
        state_var_NS = main_C_66;
      end
      main_C_66 : begin
        fsm_output = 9'b001000010;
        state_var_NS = main_C_67;
      end
      main_C_67 : begin
        fsm_output = 9'b001000011;
        state_var_NS = main_C_68;
      end
      main_C_68 : begin
        fsm_output = 9'b001000100;
        state_var_NS = main_C_69;
      end
      main_C_69 : begin
        fsm_output = 9'b001000101;
        state_var_NS = main_C_70;
      end
      main_C_70 : begin
        fsm_output = 9'b001000110;
        state_var_NS = main_C_71;
      end
      main_C_71 : begin
        fsm_output = 9'b001000111;
        state_var_NS = main_C_72;
      end
      main_C_72 : begin
        fsm_output = 9'b001001000;
        state_var_NS = main_C_73;
      end
      main_C_73 : begin
        fsm_output = 9'b001001001;
        state_var_NS = main_C_74;
      end
      main_C_74 : begin
        fsm_output = 9'b001001010;
        state_var_NS = main_C_75;
      end
      main_C_75 : begin
        fsm_output = 9'b001001011;
        state_var_NS = main_C_76;
      end
      main_C_76 : begin
        fsm_output = 9'b001001100;
        state_var_NS = main_C_77;
      end
      main_C_77 : begin
        fsm_output = 9'b001001101;
        state_var_NS = main_C_78;
      end
      main_C_78 : begin
        fsm_output = 9'b001001110;
        state_var_NS = main_C_79;
      end
      main_C_79 : begin
        fsm_output = 9'b001001111;
        state_var_NS = main_C_80;
      end
      main_C_80 : begin
        fsm_output = 9'b001010000;
        state_var_NS = main_C_81;
      end
      main_C_81 : begin
        fsm_output = 9'b001010001;
        state_var_NS = main_C_82;
      end
      main_C_82 : begin
        fsm_output = 9'b001010010;
        state_var_NS = main_C_83;
      end
      main_C_83 : begin
        fsm_output = 9'b001010011;
        state_var_NS = main_C_84;
      end
      main_C_84 : begin
        fsm_output = 9'b001010100;
        state_var_NS = main_C_85;
      end
      main_C_85 : begin
        fsm_output = 9'b001010101;
        state_var_NS = main_C_86;
      end
      main_C_86 : begin
        fsm_output = 9'b001010110;
        state_var_NS = main_C_87;
      end
      main_C_87 : begin
        fsm_output = 9'b001010111;
        state_var_NS = main_C_88;
      end
      main_C_88 : begin
        fsm_output = 9'b001011000;
        state_var_NS = main_C_89;
      end
      main_C_89 : begin
        fsm_output = 9'b001011001;
        state_var_NS = main_C_90;
      end
      main_C_90 : begin
        fsm_output = 9'b001011010;
        state_var_NS = main_C_91;
      end
      main_C_91 : begin
        fsm_output = 9'b001011011;
        state_var_NS = main_C_92;
      end
      main_C_92 : begin
        fsm_output = 9'b001011100;
        state_var_NS = main_C_93;
      end
      main_C_93 : begin
        fsm_output = 9'b001011101;
        state_var_NS = main_C_94;
      end
      main_C_94 : begin
        fsm_output = 9'b001011110;
        state_var_NS = main_C_95;
      end
      main_C_95 : begin
        fsm_output = 9'b001011111;
        state_var_NS = main_C_96;
      end
      main_C_96 : begin
        fsm_output = 9'b001100000;
        state_var_NS = main_C_97;
      end
      main_C_97 : begin
        fsm_output = 9'b001100001;
        state_var_NS = main_C_98;
      end
      main_C_98 : begin
        fsm_output = 9'b001100010;
        state_var_NS = main_C_99;
      end
      main_C_99 : begin
        fsm_output = 9'b001100011;
        state_var_NS = main_C_100;
      end
      main_C_100 : begin
        fsm_output = 9'b001100100;
        state_var_NS = main_C_101;
      end
      main_C_101 : begin
        fsm_output = 9'b001100101;
        state_var_NS = main_C_102;
      end
      main_C_102 : begin
        fsm_output = 9'b001100110;
        state_var_NS = main_C_103;
      end
      main_C_103 : begin
        fsm_output = 9'b001100111;
        state_var_NS = main_C_104;
      end
      main_C_104 : begin
        fsm_output = 9'b001101000;
        state_var_NS = main_C_105;
      end
      main_C_105 : begin
        fsm_output = 9'b001101001;
        state_var_NS = main_C_106;
      end
      main_C_106 : begin
        fsm_output = 9'b001101010;
        state_var_NS = main_C_107;
      end
      main_C_107 : begin
        fsm_output = 9'b001101011;
        state_var_NS = main_C_108;
      end
      main_C_108 : begin
        fsm_output = 9'b001101100;
        state_var_NS = main_C_109;
      end
      main_C_109 : begin
        fsm_output = 9'b001101101;
        state_var_NS = main_C_110;
      end
      main_C_110 : begin
        fsm_output = 9'b001101110;
        state_var_NS = main_C_111;
      end
      main_C_111 : begin
        fsm_output = 9'b001101111;
        state_var_NS = main_C_112;
      end
      main_C_112 : begin
        fsm_output = 9'b001110000;
        state_var_NS = main_C_113;
      end
      main_C_113 : begin
        fsm_output = 9'b001110001;
        state_var_NS = main_C_114;
      end
      main_C_114 : begin
        fsm_output = 9'b001110010;
        state_var_NS = main_C_115;
      end
      main_C_115 : begin
        fsm_output = 9'b001110011;
        state_var_NS = main_C_116;
      end
      main_C_116 : begin
        fsm_output = 9'b001110100;
        state_var_NS = main_C_117;
      end
      main_C_117 : begin
        fsm_output = 9'b001110101;
        state_var_NS = main_C_118;
      end
      main_C_118 : begin
        fsm_output = 9'b001110110;
        state_var_NS = main_C_119;
      end
      main_C_119 : begin
        fsm_output = 9'b001110111;
        state_var_NS = main_C_120;
      end
      main_C_120 : begin
        fsm_output = 9'b001111000;
        state_var_NS = main_C_121;
      end
      main_C_121 : begin
        fsm_output = 9'b001111001;
        state_var_NS = main_C_122;
      end
      main_C_122 : begin
        fsm_output = 9'b001111010;
        state_var_NS = main_C_123;
      end
      main_C_123 : begin
        fsm_output = 9'b001111011;
        state_var_NS = main_C_124;
      end
      main_C_124 : begin
        fsm_output = 9'b001111100;
        state_var_NS = main_C_125;
      end
      main_C_125 : begin
        fsm_output = 9'b001111101;
        state_var_NS = main_C_126;
      end
      main_C_126 : begin
        fsm_output = 9'b001111110;
        state_var_NS = main_C_127;
      end
      main_C_127 : begin
        fsm_output = 9'b001111111;
        state_var_NS = main_C_128;
      end
      main_C_128 : begin
        fsm_output = 9'b010000000;
        state_var_NS = main_C_129;
      end
      main_C_129 : begin
        fsm_output = 9'b010000001;
        state_var_NS = main_C_130;
      end
      main_C_130 : begin
        fsm_output = 9'b010000010;
        state_var_NS = main_C_131;
      end
      main_C_131 : begin
        fsm_output = 9'b010000011;
        state_var_NS = main_C_132;
      end
      main_C_132 : begin
        fsm_output = 9'b010000100;
        state_var_NS = main_C_133;
      end
      main_C_133 : begin
        fsm_output = 9'b010000101;
        state_var_NS = main_C_134;
      end
      main_C_134 : begin
        fsm_output = 9'b010000110;
        state_var_NS = main_C_135;
      end
      main_C_135 : begin
        fsm_output = 9'b010000111;
        state_var_NS = main_C_136;
      end
      main_C_136 : begin
        fsm_output = 9'b010001000;
        state_var_NS = main_C_137;
      end
      main_C_137 : begin
        fsm_output = 9'b010001001;
        state_var_NS = main_C_138;
      end
      main_C_138 : begin
        fsm_output = 9'b010001010;
        state_var_NS = main_C_139;
      end
      main_C_139 : begin
        fsm_output = 9'b010001011;
        state_var_NS = main_C_140;
      end
      main_C_140 : begin
        fsm_output = 9'b010001100;
        state_var_NS = main_C_141;
      end
      main_C_141 : begin
        fsm_output = 9'b010001101;
        state_var_NS = main_C_142;
      end
      main_C_142 : begin
        fsm_output = 9'b010001110;
        state_var_NS = main_C_143;
      end
      main_C_143 : begin
        fsm_output = 9'b010001111;
        state_var_NS = main_C_144;
      end
      main_C_144 : begin
        fsm_output = 9'b010010000;
        state_var_NS = main_C_145;
      end
      main_C_145 : begin
        fsm_output = 9'b010010001;
        state_var_NS = main_C_146;
      end
      main_C_146 : begin
        fsm_output = 9'b010010010;
        state_var_NS = main_C_147;
      end
      main_C_147 : begin
        fsm_output = 9'b010010011;
        state_var_NS = main_C_148;
      end
      main_C_148 : begin
        fsm_output = 9'b010010100;
        state_var_NS = main_C_149;
      end
      main_C_149 : begin
        fsm_output = 9'b010010101;
        state_var_NS = main_C_150;
      end
      main_C_150 : begin
        fsm_output = 9'b010010110;
        state_var_NS = main_C_151;
      end
      main_C_151 : begin
        fsm_output = 9'b010010111;
        state_var_NS = main_C_152;
      end
      main_C_152 : begin
        fsm_output = 9'b010011000;
        state_var_NS = main_C_153;
      end
      main_C_153 : begin
        fsm_output = 9'b010011001;
        state_var_NS = main_C_154;
      end
      main_C_154 : begin
        fsm_output = 9'b010011010;
        state_var_NS = main_C_155;
      end
      main_C_155 : begin
        fsm_output = 9'b010011011;
        state_var_NS = main_C_156;
      end
      main_C_156 : begin
        fsm_output = 9'b010011100;
        state_var_NS = main_C_157;
      end
      main_C_157 : begin
        fsm_output = 9'b010011101;
        state_var_NS = main_C_158;
      end
      main_C_158 : begin
        fsm_output = 9'b010011110;
        state_var_NS = main_C_159;
      end
      main_C_159 : begin
        fsm_output = 9'b010011111;
        state_var_NS = main_C_160;
      end
      main_C_160 : begin
        fsm_output = 9'b010100000;
        state_var_NS = main_C_161;
      end
      main_C_161 : begin
        fsm_output = 9'b010100001;
        state_var_NS = main_C_162;
      end
      main_C_162 : begin
        fsm_output = 9'b010100010;
        state_var_NS = main_C_163;
      end
      main_C_163 : begin
        fsm_output = 9'b010100011;
        state_var_NS = main_C_164;
      end
      main_C_164 : begin
        fsm_output = 9'b010100100;
        state_var_NS = main_C_165;
      end
      main_C_165 : begin
        fsm_output = 9'b010100101;
        state_var_NS = main_C_166;
      end
      main_C_166 : begin
        fsm_output = 9'b010100110;
        state_var_NS = main_C_167;
      end
      main_C_167 : begin
        fsm_output = 9'b010100111;
        state_var_NS = main_C_168;
      end
      main_C_168 : begin
        fsm_output = 9'b010101000;
        state_var_NS = main_C_169;
      end
      main_C_169 : begin
        fsm_output = 9'b010101001;
        state_var_NS = main_C_170;
      end
      main_C_170 : begin
        fsm_output = 9'b010101010;
        state_var_NS = main_C_171;
      end
      main_C_171 : begin
        fsm_output = 9'b010101011;
        state_var_NS = main_C_172;
      end
      main_C_172 : begin
        fsm_output = 9'b010101100;
        state_var_NS = main_C_173;
      end
      main_C_173 : begin
        fsm_output = 9'b010101101;
        state_var_NS = main_C_174;
      end
      main_C_174 : begin
        fsm_output = 9'b010101110;
        state_var_NS = main_C_175;
      end
      main_C_175 : begin
        fsm_output = 9'b010101111;
        state_var_NS = main_C_176;
      end
      main_C_176 : begin
        fsm_output = 9'b010110000;
        state_var_NS = main_C_177;
      end
      main_C_177 : begin
        fsm_output = 9'b010110001;
        state_var_NS = main_C_178;
      end
      main_C_178 : begin
        fsm_output = 9'b010110010;
        state_var_NS = main_C_179;
      end
      main_C_179 : begin
        fsm_output = 9'b010110011;
        state_var_NS = main_C_180;
      end
      main_C_180 : begin
        fsm_output = 9'b010110100;
        state_var_NS = main_C_181;
      end
      main_C_181 : begin
        fsm_output = 9'b010110101;
        state_var_NS = main_C_182;
      end
      main_C_182 : begin
        fsm_output = 9'b010110110;
        state_var_NS = main_C_183;
      end
      main_C_183 : begin
        fsm_output = 9'b010110111;
        state_var_NS = main_C_184;
      end
      main_C_184 : begin
        fsm_output = 9'b010111000;
        state_var_NS = main_C_185;
      end
      main_C_185 : begin
        fsm_output = 9'b010111001;
        state_var_NS = main_C_186;
      end
      main_C_186 : begin
        fsm_output = 9'b010111010;
        state_var_NS = main_C_187;
      end
      main_C_187 : begin
        fsm_output = 9'b010111011;
        state_var_NS = main_C_188;
      end
      main_C_188 : begin
        fsm_output = 9'b010111100;
        state_var_NS = main_C_189;
      end
      main_C_189 : begin
        fsm_output = 9'b010111101;
        state_var_NS = main_C_190;
      end
      main_C_190 : begin
        fsm_output = 9'b010111110;
        state_var_NS = main_C_191;
      end
      main_C_191 : begin
        fsm_output = 9'b010111111;
        state_var_NS = main_C_192;
      end
      main_C_192 : begin
        fsm_output = 9'b011000000;
        state_var_NS = main_C_193;
      end
      main_C_193 : begin
        fsm_output = 9'b011000001;
        state_var_NS = main_C_194;
      end
      main_C_194 : begin
        fsm_output = 9'b011000010;
        state_var_NS = main_C_195;
      end
      main_C_195 : begin
        fsm_output = 9'b011000011;
        state_var_NS = main_C_196;
      end
      main_C_196 : begin
        fsm_output = 9'b011000100;
        state_var_NS = main_C_197;
      end
      main_C_197 : begin
        fsm_output = 9'b011000101;
        state_var_NS = main_C_198;
      end
      main_C_198 : begin
        fsm_output = 9'b011000110;
        state_var_NS = main_C_199;
      end
      main_C_199 : begin
        fsm_output = 9'b011000111;
        state_var_NS = main_C_200;
      end
      main_C_200 : begin
        fsm_output = 9'b011001000;
        state_var_NS = main_C_201;
      end
      main_C_201 : begin
        fsm_output = 9'b011001001;
        state_var_NS = main_C_202;
      end
      main_C_202 : begin
        fsm_output = 9'b011001010;
        state_var_NS = main_C_203;
      end
      main_C_203 : begin
        fsm_output = 9'b011001011;
        state_var_NS = main_C_204;
      end
      main_C_204 : begin
        fsm_output = 9'b011001100;
        state_var_NS = main_C_205;
      end
      main_C_205 : begin
        fsm_output = 9'b011001101;
        state_var_NS = main_C_206;
      end
      main_C_206 : begin
        fsm_output = 9'b011001110;
        state_var_NS = main_C_207;
      end
      main_C_207 : begin
        fsm_output = 9'b011001111;
        state_var_NS = main_C_208;
      end
      main_C_208 : begin
        fsm_output = 9'b011010000;
        state_var_NS = main_C_209;
      end
      main_C_209 : begin
        fsm_output = 9'b011010001;
        state_var_NS = main_C_210;
      end
      main_C_210 : begin
        fsm_output = 9'b011010010;
        state_var_NS = main_C_211;
      end
      main_C_211 : begin
        fsm_output = 9'b011010011;
        state_var_NS = main_C_212;
      end
      main_C_212 : begin
        fsm_output = 9'b011010100;
        state_var_NS = main_C_213;
      end
      main_C_213 : begin
        fsm_output = 9'b011010101;
        state_var_NS = main_C_214;
      end
      main_C_214 : begin
        fsm_output = 9'b011010110;
        state_var_NS = main_C_215;
      end
      main_C_215 : begin
        fsm_output = 9'b011010111;
        state_var_NS = main_C_216;
      end
      main_C_216 : begin
        fsm_output = 9'b011011000;
        state_var_NS = main_C_217;
      end
      main_C_217 : begin
        fsm_output = 9'b011011001;
        state_var_NS = main_C_218;
      end
      main_C_218 : begin
        fsm_output = 9'b011011010;
        state_var_NS = main_C_219;
      end
      main_C_219 : begin
        fsm_output = 9'b011011011;
        state_var_NS = main_C_220;
      end
      main_C_220 : begin
        fsm_output = 9'b011011100;
        state_var_NS = main_C_221;
      end
      main_C_221 : begin
        fsm_output = 9'b011011101;
        state_var_NS = main_C_222;
      end
      main_C_222 : begin
        fsm_output = 9'b011011110;
        state_var_NS = main_C_223;
      end
      main_C_223 : begin
        fsm_output = 9'b011011111;
        state_var_NS = main_C_224;
      end
      main_C_224 : begin
        fsm_output = 9'b011100000;
        state_var_NS = main_C_225;
      end
      main_C_225 : begin
        fsm_output = 9'b011100001;
        state_var_NS = main_C_226;
      end
      main_C_226 : begin
        fsm_output = 9'b011100010;
        state_var_NS = main_C_227;
      end
      main_C_227 : begin
        fsm_output = 9'b011100011;
        state_var_NS = main_C_228;
      end
      main_C_228 : begin
        fsm_output = 9'b011100100;
        state_var_NS = main_C_229;
      end
      main_C_229 : begin
        fsm_output = 9'b011100101;
        state_var_NS = main_C_230;
      end
      main_C_230 : begin
        fsm_output = 9'b011100110;
        state_var_NS = main_C_231;
      end
      main_C_231 : begin
        fsm_output = 9'b011100111;
        state_var_NS = main_C_232;
      end
      main_C_232 : begin
        fsm_output = 9'b011101000;
        state_var_NS = main_C_233;
      end
      main_C_233 : begin
        fsm_output = 9'b011101001;
        state_var_NS = main_C_234;
      end
      main_C_234 : begin
        fsm_output = 9'b011101010;
        state_var_NS = main_C_235;
      end
      main_C_235 : begin
        fsm_output = 9'b011101011;
        state_var_NS = main_C_236;
      end
      main_C_236 : begin
        fsm_output = 9'b011101100;
        state_var_NS = main_C_237;
      end
      main_C_237 : begin
        fsm_output = 9'b011101101;
        state_var_NS = main_C_238;
      end
      main_C_238 : begin
        fsm_output = 9'b011101110;
        state_var_NS = main_C_239;
      end
      main_C_239 : begin
        fsm_output = 9'b011101111;
        state_var_NS = main_C_240;
      end
      main_C_240 : begin
        fsm_output = 9'b011110000;
        state_var_NS = main_C_241;
      end
      main_C_241 : begin
        fsm_output = 9'b011110001;
        state_var_NS = main_C_242;
      end
      main_C_242 : begin
        fsm_output = 9'b011110010;
        state_var_NS = main_C_243;
      end
      main_C_243 : begin
        fsm_output = 9'b011110011;
        state_var_NS = main_C_244;
      end
      main_C_244 : begin
        fsm_output = 9'b011110100;
        state_var_NS = main_C_245;
      end
      main_C_245 : begin
        fsm_output = 9'b011110101;
        state_var_NS = main_C_246;
      end
      main_C_246 : begin
        fsm_output = 9'b011110110;
        state_var_NS = main_C_247;
      end
      main_C_247 : begin
        fsm_output = 9'b011110111;
        state_var_NS = main_C_248;
      end
      main_C_248 : begin
        fsm_output = 9'b011111000;
        state_var_NS = main_C_249;
      end
      main_C_249 : begin
        fsm_output = 9'b011111001;
        state_var_NS = main_C_250;
      end
      main_C_250 : begin
        fsm_output = 9'b011111010;
        state_var_NS = main_C_251;
      end
      main_C_251 : begin
        fsm_output = 9'b011111011;
        state_var_NS = main_C_252;
      end
      main_C_252 : begin
        fsm_output = 9'b011111100;
        state_var_NS = main_C_253;
      end
      main_C_253 : begin
        fsm_output = 9'b011111101;
        state_var_NS = main_C_254;
      end
      main_C_254 : begin
        fsm_output = 9'b011111110;
        state_var_NS = main_C_255;
      end
      main_C_255 : begin
        fsm_output = 9'b011111111;
        state_var_NS = main_C_256;
      end
      main_C_256 : begin
        fsm_output = 9'b100000000;
        state_var_NS = main_C_257;
      end
      main_C_257 : begin
        fsm_output = 9'b100000001;
        state_var_NS = main_C_258;
      end
      main_C_258 : begin
        fsm_output = 9'b100000010;
        state_var_NS = main_C_0;
      end
      // main_C_0
      default : begin
        fsm_output = 9'b000000000;
        state_var_NS = main_C_1;
      end
    endcase
  end

  always @(posedge clk) begin
    if ( rst ) begin
      state_var <= main_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core_wait_dp
// ------------------------------------------------------------------


module fir_core_wait_dp (
  clk, rst, MAC_1_leading_sign_18_1_1_0_cmp_all_same, MAC_1_leading_sign_18_1_1_0_cmp_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same, MAC_1_leading_sign_18_1_1_0_cmp_32_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same, MAC_1_leading_sign_18_1_1_0_cmp_33_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same, MAC_1_leading_sign_18_1_1_0_cmp_34_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same, MAC_1_leading_sign_18_1_1_0_cmp_35_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same, MAC_1_leading_sign_18_1_1_0_cmp_36_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same, MAC_1_leading_sign_18_1_1_0_cmp_37_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same, MAC_1_leading_sign_18_1_1_0_cmp_38_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same, MAC_1_leading_sign_18_1_1_0_cmp_39_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same, MAC_1_leading_sign_18_1_1_0_cmp_40_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same, MAC_1_leading_sign_18_1_1_0_cmp_41_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same, MAC_1_leading_sign_18_1_1_0_cmp_42_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same, MAC_1_leading_sign_18_1_1_0_cmp_43_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same, MAC_1_leading_sign_18_1_1_0_cmp_44_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same, MAC_1_leading_sign_18_1_1_0_cmp_45_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same, MAC_1_leading_sign_18_1_1_0_cmp_46_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same, MAC_1_leading_sign_18_1_1_0_cmp_47_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same, MAC_1_leading_sign_18_1_1_0_cmp_48_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same, MAC_1_leading_sign_18_1_1_0_cmp_49_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same, MAC_1_leading_sign_18_1_1_0_cmp_50_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same, MAC_1_leading_sign_18_1_1_0_cmp_51_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same, MAC_1_leading_sign_18_1_1_0_cmp_52_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same, MAC_1_leading_sign_18_1_1_0_cmp_53_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same, MAC_1_leading_sign_18_1_1_0_cmp_54_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same, MAC_1_leading_sign_18_1_1_0_cmp_55_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same, MAC_1_leading_sign_18_1_1_0_cmp_56_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same, MAC_1_leading_sign_18_1_1_0_cmp_57_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same, MAC_1_leading_sign_18_1_1_0_cmp_58_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same, MAC_1_leading_sign_18_1_1_0_cmp_59_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same, MAC_1_leading_sign_18_1_1_0_cmp_60_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same, MAC_1_leading_sign_18_1_1_0_cmp_61_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same, MAC_1_leading_sign_18_1_1_0_cmp_62_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same, MAC_1_leading_sign_18_1_1_0_cmp_63_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg,
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg, MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg
);
  input clk;
  input rst;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  input MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;
  output MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  output MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg;
  output [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;
  reg [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;


  // Interconnect Declarations
  reg MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg;
  reg MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg;


  // Interconnect Declarations for Component Instantiations 
  assign MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg;
  assign MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg = ~ MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg;
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg <= 5'b00000;
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg <= 5'b00000;
    end
    else begin
      MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
      MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg_rneg <= ~ MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
      MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg <= MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir_core
// ------------------------------------------------------------------


module fir_core (
  clk, rst, input_m_rsc_dat, input_m_triosy_lz, input_e_rsc_dat, input_e_triosy_lz,
      taps_m_rsc_dat, taps_m_triosy_lz, taps_e_rsc_dat, taps_e_triosy_lz, return_m_rsc_dat,
      return_m_triosy_lz, return_e_rsc_dat, return_e_triosy_lz, MAC_1_leading_sign_18_1_1_0_cmp_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_all_same, MAC_1_leading_sign_18_1_1_0_cmp_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_1_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_1_rtn, MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_2_all_same, MAC_1_leading_sign_18_1_1_0_cmp_2_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_3_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_3_rtn, MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_4_all_same, MAC_1_leading_sign_18_1_1_0_cmp_4_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_5_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_5_rtn, MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_6_all_same, MAC_1_leading_sign_18_1_1_0_cmp_6_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_7_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_7_rtn, MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_8_all_same, MAC_1_leading_sign_18_1_1_0_cmp_8_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_9_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_9_rtn, MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_10_all_same, MAC_1_leading_sign_18_1_1_0_cmp_10_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_11_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_11_rtn, MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_12_all_same, MAC_1_leading_sign_18_1_1_0_cmp_12_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_13_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_13_rtn, MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_14_all_same, MAC_1_leading_sign_18_1_1_0_cmp_14_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_15_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_15_rtn, MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_16_all_same, MAC_1_leading_sign_18_1_1_0_cmp_16_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_17_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_17_rtn, MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_18_all_same, MAC_1_leading_sign_18_1_1_0_cmp_18_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_19_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_19_rtn, MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_20_all_same, MAC_1_leading_sign_18_1_1_0_cmp_20_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_21_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_21_rtn, MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_22_all_same, MAC_1_leading_sign_18_1_1_0_cmp_22_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_23_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_23_rtn, MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_24_all_same, MAC_1_leading_sign_18_1_1_0_cmp_24_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_25_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_25_rtn, MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_26_all_same, MAC_1_leading_sign_18_1_1_0_cmp_26_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_27_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_27_rtn, MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_28_all_same, MAC_1_leading_sign_18_1_1_0_cmp_28_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_29_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_29_rtn, MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_30_all_same, MAC_1_leading_sign_18_1_1_0_cmp_30_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_31_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_31_rtn, MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_32_all_same, MAC_1_leading_sign_18_1_1_0_cmp_32_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_33_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_33_rtn, MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_34_all_same, MAC_1_leading_sign_18_1_1_0_cmp_34_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_35_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_35_rtn, MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_36_all_same, MAC_1_leading_sign_18_1_1_0_cmp_36_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_37_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_37_rtn, MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_38_all_same, MAC_1_leading_sign_18_1_1_0_cmp_38_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_39_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_39_rtn, MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_40_all_same, MAC_1_leading_sign_18_1_1_0_cmp_40_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_41_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_41_rtn, MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_42_all_same, MAC_1_leading_sign_18_1_1_0_cmp_42_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_43_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_43_rtn, MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_44_all_same, MAC_1_leading_sign_18_1_1_0_cmp_44_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_45_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_45_rtn, MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_46_all_same, MAC_1_leading_sign_18_1_1_0_cmp_46_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_47_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_47_rtn, MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_48_all_same, MAC_1_leading_sign_18_1_1_0_cmp_48_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_49_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_49_rtn, MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_50_all_same, MAC_1_leading_sign_18_1_1_0_cmp_50_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_51_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_51_rtn, MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_52_all_same, MAC_1_leading_sign_18_1_1_0_cmp_52_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_53_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_53_rtn, MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_54_all_same, MAC_1_leading_sign_18_1_1_0_cmp_54_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_55_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_55_rtn, MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_56_all_same, MAC_1_leading_sign_18_1_1_0_cmp_56_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_57_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_57_rtn, MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_58_all_same, MAC_1_leading_sign_18_1_1_0_cmp_58_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_59_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_59_rtn, MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_60_all_same, MAC_1_leading_sign_18_1_1_0_cmp_60_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_61_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_61_rtn, MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa,
      MAC_1_leading_sign_18_1_1_0_cmp_62_all_same, MAC_1_leading_sign_18_1_1_0_cmp_62_rtn,
      MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa, MAC_1_leading_sign_18_1_1_0_cmp_63_all_same,
      MAC_1_leading_sign_18_1_1_0_cmp_63_rtn
);
  input clk;
  input rst;
  input [10:0] input_m_rsc_dat;
  output input_m_triosy_lz;
  input [4:0] input_e_rsc_dat;
  output input_e_triosy_lz;
  input [703:0] taps_m_rsc_dat;
  output taps_m_triosy_lz;
  input [319:0] taps_e_rsc_dat;
  output taps_e_triosy_lz;
  output [10:0] return_m_rsc_dat;
  output return_m_triosy_lz;
  output [4:0] return_e_rsc_dat;
  output return_e_triosy_lz;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  output [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  reg [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  input MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  input [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;


  // Interconnect Declarations
  wire [10:0] input_m_rsci_idat;
  wire [4:0] input_e_rsci_idat;
  wire [703:0] taps_m_rsci_idat;
  wire [319:0] taps_e_rsci_idat;
  reg [10:0] return_m_rsci_idat;
  reg [4:0] return_e_rsci_idat;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg;
  wire MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg;
  wire [8:0] fsm_output;
  wire [5:0] MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [5:0] MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire MAC_3_result_operator_result_operator_nor_tmp;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp;
  wire [5:0] MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp;
  wire [2:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp;
  wire [2:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [2:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire [3:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp;
  wire and_dcpl_1;
  wire and_dcpl_2;
  wire nor_tmp;
  wire or_tmp_6;
  wire and_dcpl_10;
  wire or_tmp_49;
  wire nor_tmp_7;
  wire mux_tmp_44;
  wire nor_tmp_10;
  wire or_tmp_116;
  wire or_dcpl_98;
  wire or_dcpl_99;
  wire or_dcpl_100;
  wire or_dcpl_103;
  wire or_dcpl_105;
  wire and_dcpl_84;
  wire and_dcpl_85;
  wire and_dcpl_86;
  wire and_dcpl_92;
  wire and_dcpl_93;
  wire and_dcpl_95;
  wire and_dcpl_97;
  wire and_dcpl_101;
  wire and_dcpl_102;
  wire and_dcpl_103;
  wire and_dcpl_105;
  wire and_dcpl_106;
  wire and_dcpl_107;
  wire and_dcpl_108;
  wire and_dcpl_109;
  wire mux_tmp_159;
  wire mux_tmp_163;
  wire or_tmp_204;
  wire nor_tmp_47;
  wire or_tmp_205;
  wire nor_tmp_49;
  wire mux_tmp_166;
  wire and_tmp_8;
  wire and_tmp_9;
  wire and_dcpl_121;
  wire mux_tmp_170;
  wire and_tmp_10;
  wire and_tmp_11;
  wire mux_tmp_172;
  wire mux_tmp_176;
  wire or_tmp_213;
  wire or_dcpl_115;
  wire nor_tmp_53;
  wire and_tmp_12;
  wire and_tmp_13;
  wire and_tmp_14;
  wire or_tmp_217;
  wire or_tmp_218;
  wire or_tmp_221;
  wire or_tmp_222;
  wire or_dcpl_120;
  wire and_dcpl_149;
  wire and_dcpl_151;
  wire and_dcpl_152;
  wire and_dcpl_153;
  wire and_dcpl_154;
  wire or_dcpl_126;
  wire and_dcpl_157;
  wire and_dcpl_158;
  wire and_dcpl_159;
  wire and_dcpl_160;
  wire and_dcpl_161;
  wire and_dcpl_162;
  wire or_dcpl_127;
  wire or_tmp_227;
  wire not_tmp_273;
  wire mux_tmp_213;
  wire mux_tmp_215;
  wire mux_tmp_217;
  wire mux_tmp_219;
  wire mux_tmp_221;
  wire mux_tmp_223;
  wire mux_tmp_225;
  wire mux_tmp_227;
  wire mux_tmp_229;
  wire and_dcpl_179;
  wire not_tmp_284;
  wire mux_tmp_232;
  wire mux_tmp_234;
  wire mux_tmp_236;
  wire mux_tmp_238;
  wire mux_tmp_240;
  wire mux_tmp_242;
  wire mux_tmp_244;
  wire and_tmp_16;
  wire and_tmp_17;
  wire and_tmp_18;
  wire and_tmp_19;
  wire and_tmp_20;
  wire and_tmp_21;
  wire and_tmp_22;
  wire or_dcpl_134;
  wire nor_tmp_66;
  wire and_dcpl_203;
  wire and_dcpl_207;
  wire and_dcpl_220;
  wire and_dcpl_221;
  wire and_dcpl_223;
  wire and_dcpl_224;
  wire and_dcpl_225;
  wire and_dcpl_235;
  wire and_dcpl_245;
  wire and_dcpl_259;
  wire and_dcpl_260;
  wire or_dcpl_150;
  wire and_dcpl_497;
  wire or_dcpl_172;
  wire mux_tmp_294;
  wire or_tmp_285;
  wire and_dcpl_546;
  wire and_dcpl_547;
  wire mux_tmp_314;
  wire or_tmp_292;
  wire or_tmp_297;
  wire or_tmp_308;
  wire or_tmp_314;
  wire or_tmp_318;
  wire or_tmp_326;
  wire or_tmp_330;
  wire or_tmp_334;
  wire or_tmp_346;
  wire or_tmp_356;
  wire or_tmp_362;
  wire or_tmp_370;
  wire or_tmp_374;
  wire and_dcpl_556;
  wire and_dcpl_561;
  wire and_dcpl_566;
  wire and_dcpl_567;
  wire and_dcpl_584;
  wire and_dcpl_585;
  wire and_dcpl_603;
  wire and_dcpl_620;
  wire and_dcpl_621;
  wire and_dcpl_626;
  wire and_dcpl_627;
  wire and_dcpl_632;
  wire and_dcpl_637;
  wire and_dcpl_690;
  wire and_dcpl_707;
  wire and_dcpl_724;
  wire and_dcpl_741;
  wire or_dcpl_278;
  wire not_tmp_640;
  wire nor_tmp_76;
  wire mux_tmp_468;
  wire or_dcpl_308;
  wire and_dcpl_910;
  wire and_dcpl_911;
  wire and_dcpl_912;
  wire and_dcpl_919;
  wire and_dcpl_921;
  wire and_dcpl_922;
  wire and_dcpl_926;
  wire and_dcpl_927;
  wire and_dcpl_928;
  wire and_dcpl_932;
  wire and_dcpl_933;
  wire and_dcpl_938;
  wire and_dcpl_939;
  wire and_dcpl_943;
  wire and_dcpl_944;
  wire and_dcpl_948;
  wire and_dcpl_949;
  wire and_dcpl_953;
  wire and_dcpl_957;
  wire and_dcpl_958;
  wire and_dcpl_962;
  wire and_dcpl_966;
  wire and_dcpl_970;
  wire and_dcpl_974;
  wire and_dcpl_981;
  wire and_dcpl_988;
  wire and_dcpl_1006;
  wire and_dcpl_1029;
  wire and_dcpl_1030;
  wire and_dcpl_1034;
  wire and_dcpl_1038;
  wire and_dcpl_1042;
  wire and_dcpl_1046;
  wire and_dcpl_1050;
  wire and_dcpl_1054;
  wire and_dcpl_1058;
  wire and_dcpl_1063;
  wire and_dcpl_1071;
  wire and_dcpl_1075;
  wire and_dcpl_1079;
  wire and_dcpl_1087;
  wire and_dcpl_1101;
  wire and_dcpl_1125;
  wire and_dcpl_1129;
  wire and_dcpl_1139;
  wire and_dcpl_1146;
  wire or_dcpl_316;
  wire mux_tmp_557;
  wire or_tmp_589;
  wire or_dcpl_368;
  wire and_dcpl_1276;
  wire and_dcpl_1287;
  wire and_dcpl_1290;
  wire and_dcpl_1291;
  wire and_dcpl_1295;
  wire and_dcpl_1298;
  wire and_dcpl_1301;
  wire and_dcpl_1304;
  wire and_dcpl_1307;
  wire and_dcpl_1326;
  wire and_dcpl_1329;
  wire and_dcpl_1332;
  wire and_dcpl_1335;
  wire and_dcpl_1338;
  wire and_dcpl_1341;
  wire and_dcpl_1344;
  wire and_dcpl_1347;
  wire and_dcpl_1427;
  wire and_dcpl_1432;
  reg ac_float_cctor_operator_return_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  reg ac_float_cctor_operator_return_9_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  reg result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  wire [10:0] MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1;
  wire MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_63_lpi_1_dfm_mx0w1;
  wire MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_62_lpi_1_dfm_mx0w1;
  wire MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_61_lpi_1_dfm_mx0w1;
  wire MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_60_lpi_1_dfm_mx0w1;
  wire MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_59_lpi_1_dfm_mx0w1;
  wire MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_58_lpi_1_dfm_mx0w1;
  wire MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_57_lpi_1_dfm_mx0w1;
  wire MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_56_lpi_1_dfm_mx0w1;
  wire MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_55_lpi_1_dfm_mx0w1;
  wire MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_54_lpi_1_dfm_mx0w1;
  wire MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_53_lpi_1_dfm_mx0w1;
  wire MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_52_lpi_1_dfm_mx0w1;
  wire MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_51_lpi_1_dfm_mx0w1;
  wire MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_50_lpi_1_dfm_mx0w1;
  wire MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_49_lpi_1_dfm_mx0w1;
  wire MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_48_lpi_1_dfm_mx0w1;
  wire MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_47_lpi_1_dfm_mx0w1;
  wire MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_46_lpi_1_dfm_mx0w1;
  wire MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_45_lpi_1_dfm_mx0w1;
  wire MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_44_lpi_1_dfm_mx0w1;
  wire MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_43_lpi_1_dfm_mx0w1;
  wire MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_42_lpi_1_dfm_mx0w1;
  wire MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_41_lpi_1_dfm_mx0w1;
  wire MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_39_lpi_1_dfm_mx0w2;
  wire MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_38_lpi_1_dfm_mx0w2;
  wire MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_37_lpi_1_dfm_mx0w2;
  wire MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_36_lpi_1_dfm_mx0w2;
  wire MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_35_lpi_1_dfm_mx0w2;
  wire MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_34_lpi_1_dfm_mx0w2;
  wire MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [10:0] MAC_ac_float_cctor_m_33_lpi_1_dfm_mx0w2;
  wire MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_33_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_32_lpi_1_dfm_mx0w2;
  wire MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_32_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w2;
  wire MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w2;
  wire MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w2;
  wire MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w2;
  wire MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w2;
  wire MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w2;
  wire MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_25_lpi_1_dfm_mx0w2;
  wire MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2;
  wire MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2;
  wire MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2;
  wire MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2;
  wire MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2;
  wire MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2;
  wire MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2;
  wire MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1;
  wire [10:0] MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w2;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva;
  reg MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva;
  reg MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva;
  reg MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva;
  reg MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva;
  reg MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva;
  reg MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva;
  reg MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva;
  reg MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva;
  reg MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva;
  reg MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva;
  reg MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva;
  reg MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva;
  reg MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva;
  reg MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva;
  reg MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva;
  reg MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva;
  reg MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva;
  reg MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva;
  reg MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva;
  reg MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva;
  reg MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva;
  reg MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva;
  reg MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva;
  reg MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva;
  reg MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva;
  reg MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva;
  reg MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva;
  reg MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva;
  reg MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva;
  reg MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva;
  reg MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva;
  reg MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva;
  reg MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva;
  reg MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva;
  reg MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva;
  reg MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva;
  reg MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva;
  reg MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva;
  reg MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva;
  reg MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva;
  reg MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva;
  reg MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva;
  reg MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva;
  reg MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva;
  reg MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva;
  reg MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva;
  reg MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva;
  reg MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva;
  reg MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva;
  reg MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva;
  reg MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva;
  reg MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva;
  reg MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva;
  reg MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva;
  reg MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva;
  reg MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva;
  reg MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva;
  reg MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva;
  reg MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva;
  reg MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva;
  reg MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva;
  reg MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva;
  reg MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1;
  wire [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1;
  reg [10:0] delay_lane_m_62_sva;
  reg [10:0] delay_lane_m_61_sva;
  reg [10:0] delay_lane_m_60_sva;
  reg [10:0] delay_lane_m_59_sva;
  reg [10:0] delay_lane_m_58_sva;
  reg [10:0] delay_lane_m_57_sva;
  reg [10:0] delay_lane_m_56_sva;
  reg [10:0] delay_lane_m_55_sva;
  reg [10:0] delay_lane_m_54_sva;
  reg [10:0] delay_lane_m_53_sva;
  reg [10:0] delay_lane_m_52_sva;
  reg [10:0] delay_lane_m_51_sva;
  reg [10:0] delay_lane_m_50_sva;
  reg [10:0] delay_lane_m_49_sva;
  reg [10:0] delay_lane_m_48_sva;
  reg [10:0] delay_lane_m_47_sva;
  reg [10:0] delay_lane_m_46_sva;
  reg [10:0] delay_lane_m_45_sva;
  reg [10:0] delay_lane_m_44_sva;
  reg [10:0] delay_lane_m_43_sva;
  reg [10:0] delay_lane_m_42_sva;
  reg [10:0] delay_lane_m_41_sva;
  reg [10:0] delay_lane_m_40_sva;
  reg [10:0] delay_lane_m_39_sva;
  reg [10:0] delay_lane_m_38_sva;
  reg [10:0] delay_lane_m_37_sva;
  reg [10:0] delay_lane_m_36_sva;
  reg [10:0] delay_lane_m_35_sva;
  reg [10:0] delay_lane_m_34_sva;
  reg [10:0] delay_lane_m_33_sva;
  reg [10:0] delay_lane_m_32_sva;
  reg [10:0] delay_lane_m_31_sva;
  reg [10:0] delay_lane_m_30_sva;
  reg [10:0] delay_lane_m_29_sva;
  reg [10:0] delay_lane_m_28_sva;
  reg [10:0] delay_lane_m_27_sva;
  reg [10:0] delay_lane_m_26_sva;
  reg [10:0] delay_lane_m_25_sva;
  reg [10:0] delay_lane_m_24_sva;
  reg [10:0] delay_lane_m_23_sva;
  reg [10:0] delay_lane_m_22_sva;
  reg [10:0] delay_lane_m_21_sva;
  reg [10:0] delay_lane_m_20_sva;
  reg [10:0] delay_lane_m_19_sva;
  reg [10:0] delay_lane_m_18_sva;
  reg [10:0] delay_lane_m_17_sva;
  reg [10:0] delay_lane_m_16_sva;
  reg [10:0] delay_lane_m_15_sva;
  reg [10:0] delay_lane_m_14_sva;
  reg [10:0] delay_lane_m_13_sva;
  reg [10:0] delay_lane_m_12_sva;
  reg [10:0] delay_lane_m_11_sva;
  reg [10:0] delay_lane_m_10_sva;
  reg [10:0] delay_lane_m_9_sva;
  reg [10:0] delay_lane_m_8_sva;
  reg [10:0] delay_lane_m_7_sva;
  reg [10:0] delay_lane_m_6_sva;
  reg [10:0] delay_lane_m_5_sva;
  reg [10:0] delay_lane_m_4_sva;
  reg [10:0] delay_lane_m_3_sva;
  reg [10:0] delay_lane_m_1_sva;
  reg [10:0] delay_lane_m_0_sva;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva;
  reg [2:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  wire [3:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva;
  reg [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_33_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_32_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0;
  wire [10:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1;
  wire [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [4:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
  wire [21:0] ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
  wire [6:0] MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_253_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_63_seb;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0;
  wire [6:0] MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_249_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_62_seb;
  wire and_221_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0;
  wire [6:0] MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_245_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_61_seb;
  wire and_220_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0;
  wire [6:0] MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_241_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_60_seb;
  wire and_219_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0;
  wire [6:0] MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_237_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_59_seb;
  wire nor_275_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0;
  wire [6:0] MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_233_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_58_seb;
  wire nor_274_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0;
  wire [6:0] MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_229_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_57_seb;
  wire nor_273_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0;
  wire [6:0] MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_225_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_56_seb;
  wire nor_272_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0;
  wire [6:0] MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_221_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_55_seb;
  wire and_210_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0;
  wire [6:0] MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_217_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_54_seb;
  wire nor_271_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0;
  wire [6:0] MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_213_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_53_seb;
  wire nor_270_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0;
  wire [6:0] MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_209_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_52_seb;
  wire nor_269_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0;
  wire [6:0] MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_205_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_51_seb;
  wire nor_268_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0;
  wire [6:0] MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_201_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_50_seb;
  wire nor_267_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0;
  wire [6:0] MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_197_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_49_seb;
  wire nor_266_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0;
  wire [6:0] MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_193_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_48_seb;
  wire nor_265_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0;
  wire [6:0] MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_189_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_47_seb;
  wire nor_264_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0;
  wire [6:0] MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_185_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_46_seb;
  wire nor_263_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0;
  wire [6:0] MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_181_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_45_seb;
  wire nor_262_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0;
  wire [6:0] MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_177_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_44_seb;
  wire and_196_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0;
  wire [6:0] MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_173_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_43_seb;
  wire nor_261_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0;
  wire [6:0] MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_169_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_42_seb;
  wire nor_260_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0;
  wire [6:0] MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_165_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_41_seb;
  wire nor_259_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0;
  wire [6:0] MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_40_seb;
  wire nor_258_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0;
  wire [6:0] MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_157_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_39_seb;
  wire nor_257_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0;
  wire [6:0] MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_153_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_38_seb;
  wire nor_256_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0;
  wire [6:0] MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_37_seb;
  wire nor_255_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0;
  wire [6:0] MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_36_seb;
  wire nor_254_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0;
  wire [6:0] MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_35_seb;
  wire nor_253_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0;
  wire [6:0] MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_34_seb;
  wire nor_252_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0;
  wire [6:0] MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [7:0] nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt;
  wire [6:0] MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire [7:0] nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_33_seb;
  wire and_184_ssc;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0;
  reg [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1;
  wire operator_13_2_true_AC_TRN_AC_WRAP_or_ssc;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse;
  wire or_741_cse;
  wire or_735_cse;
  wire nor_434_cse;
  wire nor_431_cse;
  wire nor_428_cse;
  wire nor_425_cse;
  wire nor_421_cse;
  wire nor_415_cse;
  wire nor_412_cse;
  wire nor_409_cse;
  wire nor_406_cse;
  wire nor_403_cse;
  wire nor_401_cse;
  wire nor_398_cse;
  wire nor_396_cse;
  wire or_627_cse;
  wire nor_68_cse;
  wire or_150_cse;
  wire nor_364_cse;
  wire or_452_cse;
  wire nor_360_cse;
  wire or_456_cse;
  wire nor_357_cse;
  wire nor_354_cse;
  wire nor_351_cse;
  wire nor_348_cse;
  wire nor_345_cse;
  wire and_1669_cse;
  wire nor_342_cse;
  wire nor_339_cse;
  wire nor_418_cse;
  wire nor_362_cse;
  wire or_458_cse;
  reg reg_return_e_triosy_obj_ld_cse;
  reg reg_taps_e_triosy_obj_ld_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse;
  wire operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse;
  wire nor_641_cse;
  wire and_1698_cse;
  wire nor_616_cse;
  wire nor_600_cse;
  wire nor_587_cse;
  wire nor_636_cse;
  wire nor_568_cse;
  wire or_918_cse;
  wire or_1164_cse;
  wire and_1725_cse;
  wire nor_555_cse;
  wire or_1162_cse;
  wire or_1161_cse;
  wire or_1160_cse;
  wire nor_632_cse;
  wire nor_533_cse;
  wire or_1159_cse;
  wire or_1158_cse;
  wire nor_628_cse;
  wire nor_624_cse;
  wire nor_620_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse;
  wire or_351_cse;
  wire nor_518_cse;
  wire nor_521_cse;
  wire nor_523_cse;
  wire nor_528_cse;
  wire nor_537_cse;
  wire nor_542_cse;
  wire nor_548_cse;
  wire nor_550_cse;
  wire nor_562_cse;
  wire nor_566_cse;
  wire nor_574_cse;
  wire nor_578_cse;
  wire nor_581_cse;
  wire nor_585_cse;
  wire nor_594_cse;
  wire nor_598_cse;
  wire nor_606_cse;
  wire nor_610_cse;
  wire nor_614_cse;
  wire nor_459_cse;
  wire nor_455_cse;
  wire nor_451_cse;
  wire nor_447_cse;
  wire nor_442_cse;
  wire nor_438_cse;
  wire or_969_cse;
  wire nor_225_cse;
  wire and_1670_cse;
  wire or_1120_cse;
  wire or_224_cse;
  wire or_151_cse;
  wire or_1113_cse;
  wire nor_221_cse;
  wire and_1685_cse;
  wire or_152_cse;
  wire nor_136_cse;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_cse;
  wire or_1133_cse;
  wire and_1673_cse;
  wire and_1731_cse;
  wire and_1695_cse;
  wire nor_369_cse;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc;
  reg [3:0] MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0;
  reg [3:0] MAC_ac_float_cctor_m_49_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0;
  reg MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5;
  wire or_1132_cse;
  wire or_1128_cse;
  wire mux_80_cse;
  wire mux_59_cse;
  wire or_123_cse;
  wire and_4_cse;
  wire mux_65_cse;
  wire or_1124_cse;
  wire or_tmp_717;
  wire or_tmp_718;
  wire or_tmp_719;
  wire or_tmp_725;
  wire or_tmp_731;
  wire or_tmp_734;
  wire mux_tmp;
  wire nor_tmp_132;
  wire mux_tmp_722;
  wire mux_tmp_723;
  wire mux_tmp_724;
  wire mux_tmp_725;
  wire mux_tmp_726;
  wire mux_tmp_727;
  wire mux_tmp_728;
  wire mux_tmp_729;
  wire mux_tmp_730;
  wire mux_tmp_731;
  wire mux_tmp_732;
  wire or_tmp_746;
  wire or_tmp_747;
  wire mux_tmp_733;
  wire or_tmp_748;
  wire or_tmp_762;
  wire mux_tmp_734;
  wire mux_tmp_735;
  wire nor_tmp_135;
  wire mux_tmp_736;
  wire mux_tmp_737;
  wire mux_tmp_739;
  wire mux_tmp_740;
  wire mux_tmp_741;
  wire mux_tmp_742;
  wire mux_tmp_743;
  wire mux_tmp_744;
  wire mux_tmp_745;
  wire mux_tmp_746;
  wire mux_tmp_747;
  wire mux_tmp_748;
  wire mux_tmp_750;
  wire or_tmp_774;
  wire mux_tmp_751;
  wire mux_tmp_752;
  wire or_tmp_776;
  wire or_tmp_777;
  wire or_tmp_783;
  wire nor_tmp_137;
  wire or_tmp_792;
  wire mux_tmp_754;
  wire or_tmp_793;
  wire or_tmp_794;
  wire mux_tmp_755;
  wire mux_tmp_757;
  wire mux_tmp_758;
  wire mux_tmp_759;
  wire mux_tmp_760;
  wire mux_tmp_761;
  wire mux_tmp_762;
  wire mux_tmp_763;
  wire mux_tmp_764;
  wire mux_tmp_765;
  wire mux_tmp_766;
  wire mux_tmp_767;
  wire mux_tmp_768;
  wire mux_tmp_770;
  wire mux_tmp_771;
  wire mux_tmp_772;
  wire mux_tmp_773;
  wire mux_tmp_774;
  wire mux_tmp_775;
  wire mux_tmp_776;
  wire mux_tmp_777;
  wire mux_tmp_779;
  wire mux_tmp_780;
  wire mux_tmp_781;
  wire mux_tmp_782;
  wire mux_tmp_783;
  wire mux_tmp_784;
  wire mux_tmp_785;
  wire mux_tmp_786;
  wire mux_tmp_787;
  wire mux_tmp_788;
  wire mux_tmp_791;
  wire mux_tmp_794;
  wire mux_tmp_795;
  wire mux_tmp_796;
  wire or_tmp_838;
  wire mux_tmp_801;
  wire mux_tmp_809;
  wire mux_tmp_810;
  wire or_tmp_863;
  wire or_tmp_864;
  wire or_tmp_866;
  wire or_tmp_876;
  wire mux_tmp_823;
  wire mux_tmp_824;
  wire mux_tmp_825;
  wire mux_tmp_826;
  wire mux_tmp_827;
  wire or_tmp_884;
  wire mux_tmp_829;
  wire mux_tmp_830;
  wire mux_tmp_831;
  wire mux_tmp_833;
  wire or_tmp_889;
  wire mux_tmp_834;
  wire mux_tmp_835;
  wire or_tmp_897;
  wire mux_tmp_837;
  wire mux_tmp_838;
  wire mux_tmp_839;
  wire mux_tmp_840;
  wire mux_tmp_841;
  wire mux_tmp_842;
  wire mux_tmp_843;
  wire mux_tmp_844;
  wire mux_tmp_845;
  wire mux_tmp_846;
  wire mux_tmp_847;
  wire mux_tmp_848;
  wire mux_tmp_850;
  wire mux_tmp_851;
  wire mux_tmp_852;
  wire mux_tmp_854;
  wire mux_tmp_855;
  wire mux_tmp_856;
  wire mux_tmp_857;
  wire mux_tmp_858;
  wire mux_tmp_859;
  wire mux_tmp_860;
  wire mux_tmp_861;
  wire mux_tmp_862;
  wire mux_tmp_863;
  wire mux_tmp_866;
  wire mux_tmp_869;
  wire mux_tmp_870;
  wire mux_tmp_871;
  wire mux_tmp_876;
  wire mux_tmp_884;
  wire mux_tmp_885;
  wire or_tmp_970;
  wire or_tmp_971;
  wire or_tmp_973;
  wire mux_tmp_902;
  wire mux_tmp_903;
  wire mux_tmp_904;
  wire mux_tmp_905;
  wire mux_tmp_906;
  wire or_tmp_988;
  wire mux_tmp_908;
  wire mux_tmp_909;
  wire mux_tmp_910;
  wire mux_tmp_912;
  wire or_tmp_993;
  wire mux_tmp_913;
  wire mux_tmp_914;
  wire or_tmp_1001;
  wire mux_tmp_916;
  wire mux_tmp_917;
  wire mux_tmp_918;
  wire mux_tmp_919;
  wire mux_tmp_920;
  wire mux_tmp_921;
  wire mux_tmp_922;
  wire mux_tmp_923;
  wire mux_tmp_924;
  wire mux_tmp_925;
  wire mux_tmp_926;
  wire mux_tmp_927;
  wire mux_tmp_929;
  wire mux_tmp_930;
  wire mux_tmp_931;
  wire mux_tmp_932;
  wire mux_tmp_933;
  wire mux_tmp_934;
  wire mux_tmp_935;
  wire mux_tmp_936;
  wire mux_tmp_937;
  wire mux_tmp_938;
  wire mux_tmp_939;
  wire mux_tmp_940;
  wire mux_tmp_941;
  wire mux_tmp_944;
  wire mux_tmp_947;
  wire mux_tmp_948;
  wire mux_tmp_949;
  wire mux_tmp_954;
  wire mux_tmp_962;
  wire mux_tmp_963;
  wire and_tmp_29;
  wire or_tmp_1062;
  wire or_tmp_1074;
  wire mux_tmp_976;
  wire mux_tmp_978;
  wire mux_tmp_979;
  wire mux_tmp_981;
  wire mux_tmp_982;
  wire mux_tmp_983;
  wire mux_tmp_984;
  wire or_tmp_1091;
  wire mux_tmp_986;
  wire mux_tmp_987;
  wire mux_tmp_988;
  wire mux_tmp_991;
  wire mux_tmp_994;
  wire mux_tmp_995;
  wire mux_tmp_996;
  wire mux_tmp_1001;
  wire mux_tmp_1009;
  wire mux_tmp_1010;
  reg [6:0] MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0;
  reg [6:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0;
  wire or_1557_tmp;
  wire and_1312_m1c;
  wire and_1317_m1c;
  wire and_1318_m1c;
  wire and_1321_m1c;
  wire and_1322_m1c;
  wire and_1325_m1c;
  wire and_1326_m1c;
  wire and_1328_m1c;
  wire and_1329_m1c;
  wire and_1331_m1c;
  wire and_1332_m1c;
  wire and_1334_m1c;
  wire and_1335_m1c;
  wire and_1337_m1c;
  wire and_1338_m1c;
  wire and_1339_m1c;
  wire and_1340_m1c;
  wire and_1341_m1c;
  wire and_1342_m1c;
  wire and_1343_m1c;
  wire and_1344_m1c;
  wire and_1345_m1c;
  wire and_1346_m1c;
  wire and_1347_m1c;
  wire and_1348_m1c;
  wire and_1349_m1c;
  wire and_1350_m1c;
  wire and_1351_m1c;
  wire and_1352_m1c;
  wire and_1353_m1c;
  wire and_1354_m1c;
  wire and_1356_m1c;
  wire and_1357_m1c;
  wire and_1359_m1c;
  wire and_1360_m1c;
  wire and_1362_m1c;
  wire and_1363_m1c;
  wire and_1365_m1c;
  wire and_1366_m1c;
  wire and_1368_m1c;
  wire and_1369_m1c;
  wire and_1371_m1c;
  wire and_1372_m1c;
  wire and_1374_m1c;
  wire and_1375_m1c;
  wire and_1377_m1c;
  wire and_1378_m1c;
  wire and_1379_m1c;
  wire and_1380_m1c;
  wire and_1381_m1c;
  wire and_1382_m1c;
  wire and_1383_m1c;
  wire and_1384_m1c;
  wire and_1385_m1c;
  wire and_1386_m1c;
  wire and_1387_m1c;
  wire and_1388_m1c;
  wire and_1389_m1c;
  wire and_1390_m1c;
  wire and_1391_m1c;
  wire and_1392_m1c;
  wire and_1393_m1c;
  wire and_1394_m1c;
  wire mux_1026_tmp;
  wire and_1766_cse;
  wire and_1781_cse;
  wire and_1775_cse;
  wire and_1786_cse;
  wire and_1793_cse;
  wire and_1815_cse;
  wire [5:0] MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [5:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire [6:0] nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm;
  wire mux_1035_itm;
  wire [6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm;
  wire [12:0] MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [12:0] MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [11:0] MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [11:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [12:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm;
  wire [21:0] MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [21:0] MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire [21:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm;
  wire [12:0] MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm;
  wire and_dcpl_1635;
  wire and_dcpl_1640;
  wire [6:0] z_out;
  wire [5:0] z_out_1;
  wire [6:0] nl_z_out_1;
  wire and_dcpl_1663;
  wire [10:0] z_out_2;
  reg [10:0] delay_lane_m_2_sva;
  reg [4:0] delay_lane_e_31_sva;
  reg [4:0] delay_lane_e_32_sva;
  reg [4:0] delay_lane_e_30_sva;
  reg [4:0] delay_lane_e_33_sva;
  reg [4:0] delay_lane_e_29_sva;
  reg [4:0] delay_lane_e_34_sva;
  reg [4:0] delay_lane_e_28_sva;
  reg [4:0] delay_lane_e_35_sva;
  reg [4:0] delay_lane_e_27_sva;
  reg [4:0] delay_lane_e_36_sva;
  reg [4:0] delay_lane_e_26_sva;
  reg [4:0] delay_lane_e_37_sva;
  reg [4:0] delay_lane_e_25_sva;
  reg [4:0] delay_lane_e_38_sva;
  reg [4:0] delay_lane_e_24_sva;
  reg [4:0] delay_lane_e_39_sva;
  reg [4:0] delay_lane_e_23_sva;
  reg [4:0] delay_lane_e_40_sva;
  reg [4:0] delay_lane_e_22_sva;
  reg [4:0] delay_lane_e_41_sva;
  reg [4:0] delay_lane_e_21_sva;
  reg [4:0] delay_lane_e_42_sva;
  reg [4:0] delay_lane_e_20_sva;
  reg [4:0] delay_lane_e_43_sva;
  reg [4:0] delay_lane_e_19_sva;
  reg [4:0] delay_lane_e_44_sva;
  reg [4:0] delay_lane_e_18_sva;
  reg [4:0] delay_lane_e_45_sva;
  reg [4:0] delay_lane_e_17_sva;
  reg [4:0] delay_lane_e_46_sva;
  reg [4:0] delay_lane_e_16_sva;
  reg [4:0] delay_lane_e_47_sva;
  reg [4:0] delay_lane_e_15_sva;
  reg [4:0] delay_lane_e_48_sva;
  reg [4:0] delay_lane_e_14_sva;
  reg [4:0] delay_lane_e_49_sva;
  reg [4:0] delay_lane_e_13_sva;
  reg [4:0] delay_lane_e_50_sva;
  reg [4:0] delay_lane_e_12_sva;
  reg [4:0] delay_lane_e_51_sva;
  reg [4:0] delay_lane_e_11_sva;
  reg [4:0] delay_lane_e_52_sva;
  reg [4:0] delay_lane_e_10_sva;
  reg [4:0] delay_lane_e_53_sva;
  reg [4:0] delay_lane_e_9_sva;
  reg [4:0] delay_lane_e_54_sva;
  reg [4:0] delay_lane_e_8_sva;
  reg [4:0] delay_lane_e_55_sva;
  reg [4:0] delay_lane_e_7_sva;
  reg [4:0] delay_lane_e_56_sva;
  reg [4:0] delay_lane_e_6_sva;
  reg [4:0] delay_lane_e_57_sva;
  reg [4:0] delay_lane_e_5_sva;
  reg [4:0] delay_lane_e_58_sva;
  reg [4:0] delay_lane_e_4_sva;
  reg [4:0] delay_lane_e_59_sva;
  reg [4:0] delay_lane_e_3_sva;
  reg [4:0] delay_lane_e_60_sva;
  reg [4:0] delay_lane_e_2_sva;
  reg [4:0] delay_lane_e_61_sva;
  reg [4:0] delay_lane_e_1_sva;
  reg [4:0] delay_lane_e_62_sva;
  reg [4:0] delay_lane_e_0_sva;
  reg [6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva;
  wire [7:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva;
  reg [1:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva;
  reg MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm;
  reg MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm;
  reg MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm;
  reg MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm;
  reg MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm;
  reg MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm;
  reg MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm;
  reg MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm;
  reg MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm;
  reg MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm;
  reg MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm;
  reg MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm;
  reg MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm;
  reg MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm;
  reg MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm;
  reg MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm;
  reg MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm;
  reg MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm;
  reg MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm;
  reg MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm;
  reg MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm;
  reg MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm;
  reg MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm;
  reg MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm;
  reg MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm;
  reg MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm;
  reg MAC_33_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg [3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm;
  reg MAC_34_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_35_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_36_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_37_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_38_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_39_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_40_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_41_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_42_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_43_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_44_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_45_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_46_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_47_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_48_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_49_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_50_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_51_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_52_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_53_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_54_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_55_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_56_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_57_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_58_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_59_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_60_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_61_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_62_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_63_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  reg MAC_64_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  wire return_e_rsci_idat_mx0c1;
  wire [5:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire [6:0] nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1;
  wire [11:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3;
  wire operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c1;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64;
  wire [10:0] MAC_ac_float_cctor_m_1_lpi_1_dfm_1;
  wire [3:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0;
  wire [3:0] result_m_1_lpi_1_dfm_1_10_7;
  reg [3:0] MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7;
  reg [6:0] MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0;
  reg [3:0] MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_41_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_42_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_43_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_44_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_45_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_46_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_47_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_48_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_50_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_51_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_52_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_53_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_54_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_55_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_56_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_57_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_58_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_59_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_60_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_61_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_62_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_63_lpi_1_dfm_10_7;
  reg [3:0] MAC_ac_float_cctor_m_lpi_1_dfm_10_7;
  reg MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5;
  reg [4:0] MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_10_7;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_54;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_56;
  wire leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_55;
  wire [3:0] leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_57;
  wire [5:0] operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0;
  wire [6:0] nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0;
  wire [6:0] operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0;
  wire [5:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0;
  wire [6:0] nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0;
  reg ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1;
  reg [4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2;
  reg operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0;
  reg [1:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1;
  reg [3:0] operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2;
  reg [7:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0;
  reg [3:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc;
  wire or_1042_ssc;
  wire [1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4;
  wire MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4;
  wire [3:0] MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0;
  wire result_m_1_lpi_1_dfm_1_6;
  wire [1:0] result_m_1_lpi_1_dfm_1_5_4;
  wire [3:0] result_m_1_lpi_1_dfm_1_3_0;
  wire [5:0] MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt;
  wire [6:0] nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt;
  reg result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_6;
  reg [1:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_5_4;
  wire and_568_ssc;
  wire and_573_ssc;
  wire and_575_ssc;
  wire and_579_ssc;
  wire and_584_ssc;
  wire and_589_ssc;
  wire and_595_ssc;
  wire and_599_ssc;
  wire and_603_ssc;
  wire and_607_ssc;
  wire and_613_ssc;
  wire and_617_ssc;
  wire and_621_ssc;
  wire and_625_ssc;
  wire and_631_ssc;
  wire and_635_ssc;
  wire and_639_ssc;
  wire and_643_ssc;
  wire and_649_ssc;
  wire and_655_ssc;
  wire and_660_ssc;
  wire and_665_ssc;
  wire and_669_ssc;
  wire and_673_ssc;
  wire and_677_ssc;
  wire and_681_ssc;
  wire and_685_ssc;
  wire and_689_ssc;
  wire and_693_ssc;
  wire and_697_ssc;
  wire and_701_ssc;
  wire and_705_ssc;
  wire and_709_ssc;
  wire and_713_ssc;
  wire and_718_ssc;
  wire and_722_ssc;
  wire and_726_ssc;
  wire and_730_ssc;
  wire and_735_ssc;
  wire and_739_ssc;
  wire and_743_ssc;
  wire and_747_ssc;
  wire and_752_ssc;
  wire and_756_ssc;
  wire and_760_ssc;
  wire and_764_ssc;
  wire and_769_ssc;
  wire and_773_ssc;
  wire and_777_ssc;
  wire and_781_ssc;
  wire and_785_ssc;
  wire and_789_ssc;
  wire and_793_ssc;
  wire and_797_ssc;
  wire and_801_ssc;
  wire and_805_ssc;
  wire and_809_ssc;
  wire and_813_ssc;
  wire and_817_ssc;
  wire and_821_ssc;
  wire and_825_ssc;
  wire and_829_ssc;
  wire and_833_ssc;
  wire and_837_ssc;
  wire and_841_ssc;
  wire and_845_ssc;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse;
  wire MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse;
  wire nor_773_cse;
  wire nor_774_cse;
  wire or_770_rgt;
  wire and_930_rgt;
  wire and_118_rgt;
  wire or_756_rgt;
  wire and_922_rgt;
  wire and_119_rgt;
  wire or_749_rgt;
  wire and_918_rgt;
  wire and_120_rgt;
  wire or_743_rgt;
  wire and_913_rgt;
  wire and_121_rgt;
  wire or_737_rgt;
  wire and_909_rgt;
  wire and_122_rgt;
  wire or_729_rgt;
  wire and_905_rgt;
  wire nor_248_rgt;
  wire or_723_rgt;
  wire and_901_rgt;
  wire and_125_rgt;
  wire or_717_rgt;
  wire and_897_rgt;
  wire and_127_rgt;
  wire or_710_rgt;
  wire and_893_rgt;
  wire and_129_rgt;
  wire or_704_rgt;
  wire and_890_rgt;
  wire and_133_rgt;
  wire or_697_rgt;
  wire and_884_rgt;
  wire and_135_rgt;
  wire or_683_rgt;
  wire and_876_rgt;
  wire and_137_rgt;
  wire or_675_rgt;
  wire and_872_rgt;
  wire and_138_rgt;
  wire or_667_rgt;
  wire and_868_rgt;
  wire and_139_rgt;
  wire or_660_rgt;
  wire and_864_rgt;
  wire and_140_rgt;
  wire or_653_rgt;
  wire and_860_rgt;
  wire and_141_rgt;
  wire or_646_rgt;
  wire and_856_rgt;
  wire and_142_rgt;
  wire or_639_rgt;
  wire and_852_rgt;
  wire and_143_rgt;
  wire or_631_rgt;
  wire and_848_rgt;
  wire and_144_rgt;
  wire or_470_rgt;
  wire and_559_rgt;
  wire and_145_rgt;
  wire or_453_rgt;
  wire and_551_rgt;
  wire and_146_rgt;
  wire or_445_rgt;
  wire and_547_rgt;
  wire and_149_rgt;
  wire or_437_rgt;
  wire and_543_rgt;
  wire and_151_rgt;
  wire or_430_rgt;
  wire and_539_rgt;
  wire and_153_rgt;
  wire or_422_rgt;
  wire and_535_rgt;
  wire and_155_rgt;
  wire or_415_rgt;
  wire and_531_rgt;
  wire and_156_rgt;
  wire or_408_rgt;
  wire and_527_rgt;
  wire and_158_rgt;
  wire or_401_rgt;
  wire and_523_rgt;
  wire and_159_rgt;
  wire or_763_rgt;
  wire and_926_rgt;
  wire and_160_rgt;
  wire or_690_rgt;
  wire and_880_rgt;
  wire and_161_rgt;
  wire or_462_rgt;
  wire and_555_rgt;
  wire and_162_rgt;
  wire ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse;
  wire mux_194_itm;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_95_itm;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  wire MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  wire MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  reg MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0;
  reg [3:0] MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1;
  wire and_1827_cse;
  wire and_1829_cse;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_97_m1c;

  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_63_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl;
  wire MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl;
  wire MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl;
  wire MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl;
  wire MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl;
  wire MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl;
  wire MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl;
  wire MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl;
  wire MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl;
  wire MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl;
  wire MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl;
  wire MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl;
  wire MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl;
  wire MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl;
  wire MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl;
  wire MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_14_nl;
  wire mux_91_nl;
  wire mux_485_nl;
  wire nor_458_nl;
  wire mux_484_nl;
  wire nor_457_nl;
  wire or_766_nl;
  wire mux_159_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl;
  wire mux_85_nl;
  wire mux_479_nl;
  wire nor_450_nl;
  wire mux_478_nl;
  wire nor_449_nl;
  wire or_752_nl;
  wire mux_161_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl;
  wire mux_476_nl;
  wire mux_475_nl;
  wire mux_474_nl;
  wire mux_473_nl;
  wire mux_472_nl;
  wire or_747_nl;
  wire nor_77_nl;
  wire and_1702_nl;
  wire mux_163_nl;
  wire nor_846_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl;
  wire mux_469_nl;
  wire nor_443_nl;
  wire mux_468_nl;
  wire mux_165_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl;
  wire mux_466_nl;
  wire nor_439_nl;
  wire mux_465_nl;
  wire mux_167_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl;
  wire mux_463_nl;
  wire nor_435_nl;
  wire mux_462_nl;
  wire nor_73_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl;
  wire mux_460_nl;
  wire nor_432_nl;
  wire mux_459_nl;
  wire nor_72_nl;
  wire mux_168_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl;
  wire mux_457_nl;
  wire nor_429_nl;
  wire mux_456_nl;
  wire mux_455_nl;
  wire or_715_nl;
  wire mux_170_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl;
  wire mux_453_nl;
  wire nor_426_nl;
  wire mux_452_nl;
  wire nor_71_nl;
  wire mux_172_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl;
  wire mux_451_nl;
  wire mux_450_nl;
  wire mux_449_nl;
  wire mux_448_nl;
  wire or_703_nl;
  wire or_702_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl;
  wire mux_444_nl;
  wire nor_422_nl;
  wire mux_443_nl;
  wire mux_442_nl;
  wire or_695_nl;
  wire mux_174_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl;
  wire mux_436_nl;
  wire nor_416_nl;
  wire mux_435_nl;
  wire or_681_nl;
  wire mux_434_nl;
  wire or_680_nl;
  wire mux_176_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl;
  wire or_177_nl;
  wire mux_432_nl;
  wire nor_413_nl;
  wire mux_431_nl;
  wire mux_430_nl;
  wire or_673_nl;
  wire mux_178_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl;
  wire mux_428_nl;
  wire nor_410_nl;
  wire mux_427_nl;
  wire mux_426_nl;
  wire or_665_nl;
  wire mux_180_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl;
  wire mux_423_nl;
  wire mux_422_nl;
  wire nor_407_nl;
  wire mux_421_nl;
  wire or_658_nl;
  wire mux_420_nl;
  wire or_657_nl;
  wire mux_182_nl;
  wire mux_181_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl;
  wire mux_417_nl;
  wire mux_416_nl;
  wire nor_404_nl;
  wire mux_415_nl;
  wire mux_414_nl;
  wire or_651_nl;
  wire mux_184_nl;
  wire mux_183_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_46_nl;
  wire mux_411_nl;
  wire mux_410_nl;
  wire mux_409_nl;
  wire or_645_nl;
  wire mux_408_nl;
  wire or_644_nl;
  wire mux_186_nl;
  wire mux_185_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_49_nl;
  wire mux_405_nl;
  wire mux_404_nl;
  wire nor_399_nl;
  wire mux_403_nl;
  wire mux_402_nl;
  wire or_637_nl;
  wire mux_188_nl;
  wire mux_187_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_52_nl;
  wire MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_15_nl;
  wire mux_399_nl;
  wire mux_398_nl;
  wire mux_397_nl;
  wire or_630_nl;
  wire mux_396_nl;
  wire or_629_nl;
  wire mux_190_nl;
  wire mux_189_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_55_nl;
  wire MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_16_nl;
  wire mux_193_nl;
  wire mux_192_nl;
  wire mux_191_nl;
  wire or_326_nl;
  wire MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_17_nl;
  wire mux_314_nl;
  wire mux_313_nl;
  wire nor_365_nl;
  wire mux_312_nl;
  wire mux_311_nl;
  wire or_468_nl;
  wire mux_196_nl;
  wire mux_195_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_58_nl;
  wire MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_18_nl;
  wire mux_303_nl;
  wire mux_302_nl;
  wire mux_301_nl;
  wire mux_300_nl;
  wire mux_299_nl;
  wire mux_298_nl;
  wire or_451_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_61_nl;
  wire MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_19_nl;
  wire mux_295_nl;
  wire nor_358_nl;
  wire mux_294_nl;
  wire or_443_nl;
  wire mux_293_nl;
  wire or_442_nl;
  wire mux_197_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_64_nl;
  wire MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_20_nl;
  wire mux_291_nl;
  wire nor_355_nl;
  wire mux_290_nl;
  wire mux_289_nl;
  wire or_435_nl;
  wire mux_198_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_67_nl;
  wire MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_21_nl;
  wire mux_287_nl;
  wire nor_352_nl;
  wire mux_286_nl;
  wire and_1700_nl;
  wire or_427_nl;
  wire mux_199_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_70_nl;
  wire MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_22_nl;
  wire mux_284_nl;
  wire nor_349_nl;
  wire mux_283_nl;
  wire mux_282_nl;
  wire or_420_nl;
  wire mux_200_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_73_nl;
  wire MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_23_nl;
  wire mux_280_nl;
  wire nor_346_nl;
  wire mux_279_nl;
  wire mux_278_nl;
  wire or_413_nl;
  wire mux_201_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_76_nl;
  wire MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_24_nl;
  wire mux_276_nl;
  wire nor_343_nl;
  wire mux_275_nl;
  wire mux_274_nl;
  wire or_406_nl;
  wire mux_202_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_79_nl;
  wire MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_25_nl;
  wire mux_272_nl;
  wire nor_340_nl;
  wire mux_271_nl;
  wire mux_270_nl;
  wire or_399_nl;
  wire mux_203_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_82_nl;
  wire MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_26_nl;
  wire MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_27_nl;
  wire MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_28_nl;
  wire mux_482_nl;
  wire nor_454_nl;
  wire mux_481_nl;
  wire nor_453_nl;
  wire or_759_nl;
  wire mux_205_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_85_nl;
  wire mux_440_nl;
  wire nor_419_nl;
  wire mux_439_nl;
  wire mux_438_nl;
  wire or_688_nl;
  wire mux_207_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_88_nl;
  wire mux_308_nl;
  wire mux_307_nl;
  wire mux_306_nl;
  wire mux_305_nl;
  wire or_460_nl;
  wire mux_209_nl;
  wire mux_208_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_91_nl;
  wire MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_29_nl;
  wire MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl;
  wire mux_1025_nl;
  wire mux_1024_nl;
  wire mux_1023_nl;
  wire mux_1022_nl;
  wire mux_1021_nl;
  wire mux_1020_nl;
  wire mux_1019_nl;
  wire mux_1018_nl;
  wire mux_1017_nl;
  wire mux_1016_nl;
  wire mux_1110_nl;
  wire mux_1015_nl;
  wire mux_1014_nl;
  wire mux_1011_nl;
  wire mux_1114_nl;
  wire mux_1010_nl;
  wire mux_1009_nl;
  wire mux_1008_nl;
  wire mux_1007_nl;
  wire mux_1006_nl;
  wire mux_1005_nl;
  wire mux_1003_nl;
  wire mux_1111_nl;
  wire mux_1002_nl;
  wire mux_1115_nl;
  wire mux_1001_nl;
  wire mux_1000_nl;
  wire mux_978_nl;
  wire mux_1116_nl;
  wire mux_976_nl;
  wire mux_975_nl;
  wire mux_974_nl;
  wire or_1507_nl;
  wire mux_973_nl;
  wire or_1506_nl;
  wire mux_972_nl;
  wire mux_971_nl;
  wire mux_970_nl;
  wire mux_969_nl;
  wire or_1505_nl;
  wire mux_968_nl;
  wire mux_967_nl;
  wire mux_964_nl;
  wire or_1502_nl;
  wire mux_963_nl;
  wire mux_962_nl;
  wire or_1501_nl;
  wire mux_961_nl;
  wire or_1500_nl;
  wire mux_960_nl;
  wire mux_959_nl;
  wire mux_958_nl;
  wire mux_956_nl;
  wire mux_955_nl;
  wire or_1498_nl;
  wire mux_954_nl;
  wire mux_953_nl;
  wire mux_918_nl;
  wire or_1563_nl;
  wire mux_1037_nl;
  wire mux_901_nl;
  wire and_1749_nl;
  wire or_1413_nl;
  wire or_nl;
  wire or_1564_nl;
  wire mux_1038_nl;
  wire mux_898_nl;
  wire mux_897_nl;
  wire mux_896_nl;
  wire or_1410_nl;
  wire mux_895_nl;
  wire or_1409_nl;
  wire mux_894_nl;
  wire mux_893_nl;
  wire mux_892_nl;
  wire mux_891_nl;
  wire or_1408_nl;
  wire mux_890_nl;
  wire mux_889_nl;
  wire mux_886_nl;
  wire or_1405_nl;
  wire mux_885_nl;
  wire mux_884_nl;
  wire or_1404_nl;
  wire mux_883_nl;
  wire or_1403_nl;
  wire mux_882_nl;
  wire mux_881_nl;
  wire mux_880_nl;
  wire mux_878_nl;
  wire mux_877_nl;
  wire or_1401_nl;
  wire mux_876_nl;
  wire mux_875_nl;
  wire mux_839_nl;
  wire mux_823_nl;
  wire mux_822_nl;
  wire mux_821_nl;
  wire or_1306_nl;
  wire mux_820_nl;
  wire or_1304_nl;
  wire mux_819_nl;
  wire mux_818_nl;
  wire mux_817_nl;
  wire mux_816_nl;
  wire or_1303_nl;
  wire mux_815_nl;
  wire mux_814_nl;
  wire mux_811_nl;
  wire or_1298_nl;
  wire mux_810_nl;
  wire mux_809_nl;
  wire or_1297_nl;
  wire mux_808_nl;
  wire or_1295_nl;
  wire mux_807_nl;
  wire mux_806_nl;
  wire mux_805_nl;
  wire mux_803_nl;
  wire mux_802_nl;
  wire or_1293_nl;
  wire mux_801_nl;
  wire mux_800_nl;
  wire mux_756_nl;
  wire MAC_10_r_ac_float_else_and_nl;
  wire[4:0] MAC_10_r_ac_float_else_and_1_nl;
  wire mux_723_nl;
  wire mux_722_nl;
  wire mux_721_nl;
  wire mux_720_nl;
  wire mux_719_nl;
  wire and_1740_nl;
  wire mux_718_nl;
  wire nor_646_nl;
  wire or_1102_nl;
  wire mux_717_nl;
  wire mux_716_nl;
  wire nor_647_nl;
  wire or_1100_nl;
  wire mux_715_nl;
  wire nor_648_nl;
  wire or_1098_nl;
  wire mux_714_nl;
  wire mux_713_nl;
  wire mux_712_nl;
  wire nor_649_nl;
  wire or_1096_nl;
  wire mux_711_nl;
  wire nor_650_nl;
  wire or_1094_nl;
  wire mux_710_nl;
  wire mux_709_nl;
  wire nor_651_nl;
  wire or_1092_nl;
  wire mux_708_nl;
  wire nor_652_nl;
  wire or_1090_nl;
  wire mux_707_nl;
  wire mux_706_nl;
  wire mux_705_nl;
  wire mux_704_nl;
  wire nor_653_nl;
  wire or_1088_nl;
  wire mux_703_nl;
  wire and_1741_nl;
  wire or_1087_nl;
  wire mux_702_nl;
  wire mux_701_nl;
  wire nor_654_nl;
  wire or_1085_nl;
  wire mux_700_nl;
  wire nor_655_nl;
  wire or_1083_nl;
  wire mux_699_nl;
  wire mux_698_nl;
  wire mux_697_nl;
  wire and_1742_nl;
  wire or_1082_nl;
  wire mux_696_nl;
  wire and_1743_nl;
  wire or_1081_nl;
  wire mux_695_nl;
  wire mux_694_nl;
  wire and_1744_nl;
  wire or_1080_nl;
  wire mux_693_nl;
  wire nor_656_nl;
  wire or_1078_nl;
  wire mux_692_nl;
  wire mux_691_nl;
  wire mux_690_nl;
  wire mux_689_nl;
  wire mux_688_nl;
  wire and_1745_nl;
  wire or_1077_nl;
  wire mux_687_nl;
  wire and_1746_nl;
  wire or_1076_nl;
  wire mux_686_nl;
  wire mux_685_nl;
  wire nor_657_nl;
  wire or_1074_nl;
  wire mux_684_nl;
  wire and_1747_nl;
  wire or_1073_nl;
  wire mux_683_nl;
  wire mux_682_nl;
  wire mux_681_nl;
  wire nor_658_nl;
  wire or_1071_nl;
  wire mux_680_nl;
  wire nor_659_nl;
  wire or_1069_nl;
  wire mux_679_nl;
  wire mux_678_nl;
  wire nor_660_nl;
  wire or_1067_nl;
  wire mux_677_nl;
  wire nor_661_nl;
  wire or_1065_nl;
  wire mux_676_nl;
  wire mux_675_nl;
  wire mux_674_nl;
  wire mux_673_nl;
  wire nor_662_nl;
  wire or_1063_nl;
  wire mux_672_nl;
  wire nor_663_nl;
  wire or_1061_nl;
  wire mux_671_nl;
  wire mux_670_nl;
  wire nor_664_nl;
  wire or_1059_nl;
  wire mux_669_nl;
  wire nor_665_nl;
  wire or_1057_nl;
  wire mux_668_nl;
  wire mux_667_nl;
  wire mux_666_nl;
  wire nor_666_nl;
  wire or_1055_nl;
  wire mux_665_nl;
  wire nor_667_nl;
  wire or_1053_nl;
  wire mux_664_nl;
  wire mux_663_nl;
  wire nor_668_nl;
  wire or_1051_nl;
  wire mux_662_nl;
  wire and_1748_nl;
  wire or_1050_nl;
  wire mux_1109_nl;
  wire nand_150_nl;
  wire mux_1108_nl;
  wire mux_1107_nl;
  wire mux_1106_nl;
  wire mux_1105_nl;
  wire mux_1104_nl;
  wire and_1933_nl;
  wire mux_1103_nl;
  wire nand_88_nl;
  wire nand_89_nl;
  wire mux_1102_nl;
  wire mux_1101_nl;
  wire nand_90_nl;
  wire nand_91_nl;
  wire mux_1100_nl;
  wire nand_92_nl;
  wire nand_93_nl;
  wire mux_1099_nl;
  wire mux_1098_nl;
  wire mux_1097_nl;
  wire nand_94_nl;
  wire nand_95_nl;
  wire mux_1096_nl;
  wire nand_96_nl;
  wire nand_97_nl;
  wire mux_1095_nl;
  wire mux_1094_nl;
  wire nand_98_nl;
  wire nand_99_nl;
  wire mux_1093_nl;
  wire nand_100_nl;
  wire nand_101_nl;
  wire mux_1092_nl;
  wire mux_1091_nl;
  wire mux_1090_nl;
  wire mux_1089_nl;
  wire nand_102_nl;
  wire nand_103_nl;
  wire mux_1088_nl;
  wire nand_104_nl;
  wire nand_105_nl;
  wire mux_1087_nl;
  wire mux_1086_nl;
  wire nand_106_nl;
  wire nand_107_nl;
  wire mux_1085_nl;
  wire nand_108_nl;
  wire nand_109_nl;
  wire mux_1084_nl;
  wire mux_1083_nl;
  wire mux_1082_nl;
  wire nand_110_nl;
  wire nand_111_nl;
  wire mux_1081_nl;
  wire nand_112_nl;
  wire nand_113_nl;
  wire mux_1080_nl;
  wire mux_1079_nl;
  wire nand_114_nl;
  wire nand_115_nl;
  wire mux_1078_nl;
  wire nand_116_nl;
  wire nand_117_nl;
  wire mux_1077_nl;
  wire mux_1076_nl;
  wire mux_1075_nl;
  wire mux_1074_nl;
  wire mux_1073_nl;
  wire nand_118_nl;
  wire nand_119_nl;
  wire mux_1072_nl;
  wire nand_120_nl;
  wire nand_121_nl;
  wire mux_1071_nl;
  wire mux_1070_nl;
  wire nand_122_nl;
  wire nand_123_nl;
  wire mux_1069_nl;
  wire nand_124_nl;
  wire nand_125_nl;
  wire mux_1068_nl;
  wire mux_1067_nl;
  wire mux_1066_nl;
  wire nand_126_nl;
  wire nand_127_nl;
  wire mux_1065_nl;
  wire nand_128_nl;
  wire nand_129_nl;
  wire mux_1064_nl;
  wire mux_1063_nl;
  wire nand_130_nl;
  wire nand_131_nl;
  wire mux_1062_nl;
  wire nand_132_nl;
  wire nand_133_nl;
  wire mux_1061_nl;
  wire mux_1060_nl;
  wire mux_1059_nl;
  wire mux_1058_nl;
  wire nand_134_nl;
  wire nand_135_nl;
  wire mux_1057_nl;
  wire nand_136_nl;
  wire nand_137_nl;
  wire mux_1056_nl;
  wire mux_1055_nl;
  wire nand_138_nl;
  wire nand_139_nl;
  wire mux_1054_nl;
  wire nand_140_nl;
  wire nand_141_nl;
  wire mux_1053_nl;
  wire mux_1052_nl;
  wire mux_1051_nl;
  wire nand_142_nl;
  wire nand_143_nl;
  wire mux_1050_nl;
  wire nand_144_nl;
  wire nand_145_nl;
  wire mux_1049_nl;
  wire mux_1048_nl;
  wire nand_146_nl;
  wire nand_147_nl;
  wire mux_1047_nl;
  wire nand_148_nl;
  wire nand_149_nl;
  wire nor_845_nl;
  wire mux_213_nl;
  wire nor_250_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_61_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_124_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_91_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_33_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_312_nl;
  wire mux_656_nl;
  wire nor_642_nl;
  wire mux_655_nl;
  wire nor_640_nl;
  wire or_1036_nl;
  wire and_1301_nl;
  wire mux_657_nl;
  wire mux_215_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_60_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_90_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_68_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_310_nl;
  wire mux_638_nl;
  wire mux_637_nl;
  wire nor_617_nl;
  wire mux_636_nl;
  wire or_995_nl;
  wire and_1733_nl;
  wire or_991_nl;
  wire and_1277_nl;
  wire mux_639_nl;
  wire mux_217_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_59_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_89_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_92_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_308_nl;
  wire mux_634_nl;
  wire nor_613_nl;
  wire mux_633_nl;
  wire nor_612_nl;
  wire and_1273_nl;
  wire mux_635_nl;
  wire mux_219_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_88_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_72_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_36_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_306_nl;
  wire mux_631_nl;
  wire nor_609_nl;
  wire mux_630_nl;
  wire nor_608_nl;
  wire and_1269_nl;
  wire mux_632_nl;
  wire mux_221_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_57_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_120_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_87_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_74_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_304_nl;
  wire mux_628_nl;
  wire nor_605_nl;
  wire mux_627_nl;
  wire nor_604_nl;
  wire and_1265_nl;
  wire mux_629_nl;
  wire mux_223_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_56_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_86_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_76_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_302_nl;
  wire mux_625_nl;
  wire mux_624_nl;
  wire mux_623_nl;
  wire nor_601_nl;
  wire mux_622_nl;
  wire or_968_nl;
  wire and_1730_nl;
  wire and_1261_nl;
  wire mux_626_nl;
  wire mux_225_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_55_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_85_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_78_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_39_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_300_nl;
  wire mux_620_nl;
  wire nor_597_nl;
  wire mux_619_nl;
  wire nor_596_nl;
  wire and_1257_nl;
  wire mux_621_nl;
  wire mux_227_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_84_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_80_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_40_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_298_nl;
  wire mux_617_nl;
  wire nor_593_nl;
  wire mux_616_nl;
  wire nor_592_nl;
  wire and_1253_nl;
  wire mux_618_nl;
  wire mux_229_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_53_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_116_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_83_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_82_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_41_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_296_nl;
  wire mux_614_nl;
  wire mux_613_nl;
  wire nor_588_nl;
  wire mux_612_nl;
  wire or_950_nl;
  wire and_1246_nl;
  wire and_1249_nl;
  wire mux_615_nl;
  wire mux_231_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_52_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_82_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_84_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_294_nl;
  wire mux_610_nl;
  wire nor_584_nl;
  wire mux_609_nl;
  wire nor_583_nl;
  wire and_1244_nl;
  wire mux_611_nl;
  wire mux_233_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_81_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_86_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_43_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_292_nl;
  wire mux_607_nl;
  wire nor_580_nl;
  wire mux_606_nl;
  wire mux_605_nl;
  wire or_935_nl;
  wire and_1237_nl;
  wire and_1240_nl;
  wire mux_608_nl;
  wire mux_234_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_80_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_88_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_44_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_291_nl;
  wire mux_653_nl;
  wire nor_638_nl;
  wire mux_652_nl;
  wire and_1738_nl;
  wire and_1297_nl;
  wire mux_654_nl;
  wire mux_236_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_79_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_90_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_45_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_289_nl;
  wire mux_603_nl;
  wire nor_577_nl;
  wire mux_602_nl;
  wire nor_576_nl;
  wire and_1235_nl;
  wire mux_604_nl;
  wire mux_238_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_48_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_78_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_92_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_287_nl;
  wire mux_600_nl;
  wire nor_573_nl;
  wire mux_599_nl;
  wire nor_572_nl;
  wire and_1231_nl;
  wire mux_601_nl;
  wire mux_240_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_47_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_77_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_94_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_285_nl;
  wire mux_597_nl;
  wire mux_596_nl;
  wire nor_569_nl;
  wire mux_595_nl;
  wire or_917_nl;
  wire and_1724_nl;
  wire and_1227_nl;
  wire mux_598_nl;
  wire mux_242_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_76_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_96_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_48_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_283_nl;
  wire mux_593_nl;
  wire nor_565_nl;
  wire mux_592_nl;
  wire nor_564_nl;
  wire and_1223_nl;
  wire mux_594_nl;
  wire mux_244_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_45_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_75_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_49_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_281_nl;
  wire mux_590_nl;
  wire nor_561_nl;
  wire mux_589_nl;
  wire nor_560_nl;
  wire and_1219_nl;
  wire mux_591_nl;
  wire mux_246_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_44_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_74_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_100_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_279_nl;
  wire mux_587_nl;
  wire mux_586_nl;
  wire nor_556_nl;
  wire mux_585_nl;
  wire or_897_nl;
  wire and_1212_nl;
  wire and_1215_nl;
  wire mux_588_nl;
  wire mux_248_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_73_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_51_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_277_nl;
  wire mux_583_nl;
  wire nor_552_nl;
  wire and_1210_nl;
  wire mux_584_nl;
  wire mux_249_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_72_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_104_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_52_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_275_nl;
  wire mux_581_nl;
  wire nor_547_nl;
  wire mux_580_nl;
  wire mux_579_nl;
  wire or_882_nl;
  wire and_1203_nl;
  wire and_1206_nl;
  wire mux_582_nl;
  wire mux_250_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_71_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_53_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_273_nl;
  wire mux_577_nl;
  wire nor_544_nl;
  wire and_1201_nl;
  wire mux_578_nl;
  wire mux_251_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_70_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_108_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_271_nl;
  wire mux_575_nl;
  wire nor_539_nl;
  wire and_1197_nl;
  wire mux_576_nl;
  wire mux_252_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_69_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_55_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_270_nl;
  wire mux_650_nl;
  wire nor_634_nl;
  wire mux_649_nl;
  wire and_1737_nl;
  wire and_1293_nl;
  wire mux_651_nl;
  wire mux_253_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_68_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_112_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_56_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_268_nl;
  wire mux_573_nl;
  wire mux_572_nl;
  wire nor_534_nl;
  wire mux_571_nl;
  wire or_864_nl;
  wire or_863_nl;
  wire and_1714_nl;
  wire and_1715_nl;
  wire and_1193_nl;
  wire mux_574_nl;
  wire mux_254_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_67_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_114_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_57_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_266_nl;
  wire mux_569_nl;
  wire nor_530_nl;
  wire and_1189_nl;
  wire mux_570_nl;
  wire mux_255_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_66_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_116_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_264_nl;
  wire mux_567_nl;
  wire nor_525_nl;
  wire and_1185_nl;
  wire mux_568_nl;
  wire mux_256_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_65_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_118_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_59_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_262_nl;
  wire mux_565_nl;
  wire mux_564_nl;
  wire nor_520_nl;
  wire mux_563_nl;
  wire mux_562_nl;
  wire mux_561_nl;
  wire or_844_nl;
  wire and_1181_nl;
  wire mux_566_nl;
  wire mux_257_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_64_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_120_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_60_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_261_nl;
  wire mux_647_nl;
  wire nor_630_nl;
  wire mux_646_nl;
  wire and_1736_nl;
  wire and_1289_nl;
  wire mux_648_nl;
  wire mux_258_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_96_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_63_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_122_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_61_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_260_nl;
  wire mux_644_nl;
  wire nor_626_nl;
  wire mux_643_nl;
  wire and_1735_nl;
  wire and_1285_nl;
  wire mux_645_nl;
  wire mux_259_nl;
  wire nor_138_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_62_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_124_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_259_nl;
  wire mux_641_nl;
  wire nor_622_nl;
  wire mux_640_nl;
  wire and_1734_nl;
  wire and_1281_nl;
  wire mux_642_nl;
  wire[2:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[3:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire MAC_3_r_ac_float_else_and_nl;
  wire[4:0] MAC_3_r_ac_float_else_and_1_nl;
  wire mux_260_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl;
  wire[1:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_64_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_126_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_63_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl;
  wire mux_261_nl;
  wire mux_559_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[1:0] MAC_11_r_ac_float_else_and_nl;
  wire[3:0] MAC_11_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_12_r_ac_float_else_and_nl;
  wire[4:0] MAC_12_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_13_r_ac_float_else_and_nl;
  wire[4:0] MAC_13_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_14_r_ac_float_else_and_nl;
  wire[4:0] MAC_14_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_15_r_ac_float_else_and_nl;
  wire[4:0] MAC_15_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_16_r_ac_float_else_and_nl;
  wire[4:0] MAC_16_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_17_r_ac_float_else_and_nl;
  wire[4:0] MAC_17_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_18_r_ac_float_else_and_nl;
  wire[4:0] MAC_18_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_19_r_ac_float_else_and_nl;
  wire[4:0] MAC_19_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_2_r_ac_float_else_and_nl;
  wire[4:0] MAC_2_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_20_r_ac_float_else_and_nl;
  wire[4:0] MAC_20_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_21_r_ac_float_else_and_nl;
  wire MAC_21_r_ac_float_else_and_1_nl;
  wire[3:0] MAC_21_r_ac_float_else_and_2_nl;
  wire[6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_22_r_ac_float_else_and_nl;
  wire[4:0] MAC_22_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_23_r_ac_float_else_and_nl;
  wire[4:0] MAC_23_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_24_r_ac_float_else_and_nl;
  wire[4:0] MAC_24_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_25_r_ac_float_else_and_nl;
  wire[4:0] MAC_25_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_26_r_ac_float_else_and_nl;
  wire[4:0] MAC_26_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_27_r_ac_float_else_and_nl;
  wire[4:0] MAC_27_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_28_r_ac_float_else_and_nl;
  wire[4:0] MAC_28_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_29_r_ac_float_else_and_nl;
  wire[4:0] MAC_29_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_30_r_ac_float_else_and_nl;
  wire[4:0] MAC_30_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_31_r_ac_float_else_and_nl;
  wire[4:0] MAC_31_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_32_r_ac_float_else_and_nl;
  wire[4:0] MAC_32_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_33_r_ac_float_else_and_nl;
  wire[4:0] MAC_33_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_4_r_ac_float_else_and_nl;
  wire[4:0] MAC_4_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_5_r_ac_float_else_and_nl;
  wire[4:0] MAC_5_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_6_r_ac_float_else_and_nl;
  wire[4:0] MAC_6_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_7_r_ac_float_else_and_nl;
  wire[4:0] MAC_7_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_8_r_ac_float_else_and_nl;
  wire[4:0] MAC_8_r_ac_float_else_and_1_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl;
  wire MAC_9_r_ac_float_else_and_nl;
  wire[4:0] MAC_9_r_ac_float_else_and_1_nl;
  wire MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire and_251_nl;
  wire and_254_nl;
  wire and_257_nl;
  wire MAC_33_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire and_261_nl;
  wire and_264_nl;
  wire and_267_nl;
  wire MAC_34_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire MAC_35_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire MAC_36_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_43_nl;
  wire and_274_nl;
  wire MAC_37_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_44_nl;
  wire and_276_nl;
  wire MAC_38_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire and_279_nl;
  wire and_284_nl;
  wire and_287_nl;
  wire MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_27_nl;
  wire and_289_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_51_nl;
  wire[3:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_28_nl;
  wire and_291_nl;
  wire MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_29_nl;
  wire and_293_nl;
  wire MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_30_nl;
  wire and_295_nl;
  wire MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_31_nl;
  wire and_297_nl;
  wire MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_32_nl;
  wire and_299_nl;
  wire MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_33_nl;
  wire and_301_nl;
  wire MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_34_nl;
  wire and_303_nl;
  wire MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_35_nl;
  wire and_305_nl;
  wire MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_36_nl;
  wire and_307_nl;
  wire MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_37_nl;
  wire and_309_nl;
  wire MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_39_nl;
  wire and_311_nl;
  wire MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_40_nl;
  wire and_313_nl;
  wire MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_298_nl;
  wire and_315_nl;
  wire MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_299_nl;
  wire and_317_nl;
  wire MAC_25_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_300_nl;
  wire and_319_nl;
  wire MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_301_nl;
  wire and_321_nl;
  wire MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_302_nl;
  wire and_323_nl;
  wire MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_303_nl;
  wire and_325_nl;
  wire MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_304_nl;
  wire and_327_nl;
  wire MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_305_nl;
  wire and_329_nl;
  wire MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_306_nl;
  wire and_331_nl;
  wire MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire[3:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire nor_307_nl;
  wire and_333_nl;
  wire MAC_32_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_nl;
  wire MAC_59_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_nl;
  wire MAC_58_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_nl;
  wire MAC_57_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_nl;
  wire MAC_55_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_nl;
  wire MAC_54_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_nl;
  wire MAC_53_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_nl;
  wire MAC_52_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_nl;
  wire MAC_51_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_nl;
  wire MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_nl;
  wire MAC_50_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_nl;
  wire MAC_49_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_nl;
  wire MAC_48_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_nl;
  wire MAC_47_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_nl;
  wire MAC_46_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_nl;
  wire MAC_45_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_nl;
  wire MAC_44_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl;
  wire MAC_43_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl;
  wire MAC_42_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl;
  wire MAC_41_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl;
  wire MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl;
  wire MAC_39_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl;
  wire MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl;
  wire MAC_63_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl;
  wire MAC_62_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl;
  wire MAC_61_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl;
  wire MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl;
  wire MAC_60_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl;
  wire MAC_56_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl;
  wire[3:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl;
  wire and_270_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[10:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_128_nl;
  wire[10:0] result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl;
  wire[1:0] MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[1:0] MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire[2:0] nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl;
  wire MAC_34_r_ac_float_else_and_nl;
  wire[4:0] MAC_34_r_ac_float_else_and_1_nl;
  wire MAC_35_r_ac_float_else_and_nl;
  wire[4:0] MAC_35_r_ac_float_else_and_1_nl;
  wire MAC_36_r_ac_float_else_and_nl;
  wire[4:0] MAC_36_r_ac_float_else_and_1_nl;
  wire MAC_37_r_ac_float_else_and_nl;
  wire[4:0] MAC_37_r_ac_float_else_and_1_nl;
  wire MAC_38_r_ac_float_else_and_nl;
  wire[4:0] MAC_38_r_ac_float_else_and_1_nl;
  wire MAC_39_r_ac_float_else_and_nl;
  wire[4:0] MAC_39_r_ac_float_else_and_1_nl;
  wire MAC_40_r_ac_float_else_and_nl;
  wire[4:0] MAC_40_r_ac_float_else_and_1_nl;
  wire MAC_41_r_ac_float_else_and_nl;
  wire[4:0] MAC_41_r_ac_float_else_and_1_nl;
  wire MAC_42_r_ac_float_else_and_nl;
  wire[4:0] MAC_42_r_ac_float_else_and_1_nl;
  wire MAC_43_r_ac_float_else_and_nl;
  wire[4:0] MAC_43_r_ac_float_else_and_1_nl;
  wire MAC_44_r_ac_float_else_and_nl;
  wire[4:0] MAC_44_r_ac_float_else_and_1_nl;
  wire MAC_45_r_ac_float_else_and_nl;
  wire[4:0] MAC_45_r_ac_float_else_and_1_nl;
  wire MAC_46_r_ac_float_else_and_nl;
  wire[4:0] MAC_46_r_ac_float_else_and_1_nl;
  wire MAC_47_r_ac_float_else_and_nl;
  wire[4:0] MAC_47_r_ac_float_else_and_1_nl;
  wire MAC_48_r_ac_float_else_and_nl;
  wire[4:0] MAC_48_r_ac_float_else_and_1_nl;
  wire MAC_49_r_ac_float_else_and_nl;
  wire[4:0] MAC_49_r_ac_float_else_and_1_nl;
  wire MAC_50_r_ac_float_else_and_nl;
  wire[4:0] MAC_50_r_ac_float_else_and_1_nl;
  wire MAC_51_r_ac_float_else_and_nl;
  wire[4:0] MAC_51_r_ac_float_else_and_1_nl;
  wire MAC_52_r_ac_float_else_and_nl;
  wire[4:0] MAC_52_r_ac_float_else_and_1_nl;
  wire MAC_53_r_ac_float_else_and_nl;
  wire[4:0] MAC_53_r_ac_float_else_and_1_nl;
  wire MAC_54_r_ac_float_else_and_nl;
  wire[4:0] MAC_54_r_ac_float_else_and_1_nl;
  wire MAC_55_r_ac_float_else_and_nl;
  wire[4:0] MAC_55_r_ac_float_else_and_1_nl;
  wire MAC_56_r_ac_float_else_and_nl;
  wire[4:0] MAC_56_r_ac_float_else_and_1_nl;
  wire MAC_57_r_ac_float_else_and_nl;
  wire[4:0] MAC_57_r_ac_float_else_and_1_nl;
  wire MAC_58_r_ac_float_else_and_nl;
  wire[4:0] MAC_58_r_ac_float_else_and_1_nl;
  wire MAC_59_r_ac_float_else_and_nl;
  wire[4:0] MAC_59_r_ac_float_else_and_1_nl;
  wire MAC_60_r_ac_float_else_and_nl;
  wire[4:0] MAC_60_r_ac_float_else_and_1_nl;
  wire MAC_61_r_ac_float_else_and_nl;
  wire[4:0] MAC_61_r_ac_float_else_and_1_nl;
  wire MAC_62_r_ac_float_else_and_nl;
  wire[4:0] MAC_62_r_ac_float_else_and_1_nl;
  wire MAC_63_r_ac_float_else_and_nl;
  wire[4:0] MAC_63_r_ac_float_else_and_1_nl;
  wire MAC_1_r_ac_float_else_and_nl;
  wire[4:0] MAC_1_r_ac_float_else_and_1_nl;
  wire MAC_64_r_ac_float_else_and_nl;
  wire[4:0] MAC_64_r_ac_float_else_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_166_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_167_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_170_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_171_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_174_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_175_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_178_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_179_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_182_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_183_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_186_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_187_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_190_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_191_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_194_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_195_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_198_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_199_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_202_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_203_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_206_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_207_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_210_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_211_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_214_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_215_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_218_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_219_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_222_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_223_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_226_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_227_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_230_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_231_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_234_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_235_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_238_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_239_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_242_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_243_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_246_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_247_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_250_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_251_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_254_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_255_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl;
  wire[6:0] MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl;
  wire[6:0] MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl;
  wire[6:0] MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl;
  wire[6:0] MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl;
  wire[6:0] MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl;
  wire[6:0] MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl;
  wire[6:0] MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl;
  wire[6:0] MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl;
  wire[6:0] MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl;
  wire[6:0] MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl;
  wire[6:0] MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl;
  wire[6:0] MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl;
  wire[6:0] MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl;
  wire[6:0] MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl;
  wire[6:0] MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl;
  wire[6:0] MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl;
  wire[6:0] MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl;
  wire[6:0] MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl;
  wire[6:0] MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl;
  wire[6:0] MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl;
  wire[6:0] MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl;
  wire[6:0] MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl;
  wire[6:0] MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_130_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl;
  wire[6:0] MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl;
  wire[6:0] MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_138_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl;
  wire[6:0] MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_142_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl;
  wire[6:0] MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_146_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl;
  wire[6:0] MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_150_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl;
  wire[6:0] MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_154_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_155_nl;
  wire[6:0] MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl;
  wire[6:0] MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_32_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_129_nl;
  wire[6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_nl;
  wire[6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl;
  wire[6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl;
  wire[6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl;
  wire[6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl;
  wire[6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl;
  wire[6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl;
  wire[6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl;
  wire[6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl;
  wire[6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl;
  wire[6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl;
  wire[6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl;
  wire[6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl;
  wire[6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl;
  wire[6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl;
  wire ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl;
  wire[5:0] MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_195_nl;
  wire[1:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_318_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_260_nl;
  wire[3:0] result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_319_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_261_nl;
  wire[6:0] MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl;
  wire[7:0] nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl;
  wire[5:0] MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire or_320_nl;
  wire mux_204_nl;
  wire mux_214_nl;
  wire and_1684_nl;
  wire or_360_nl;
  wire or_361_nl;
  wire or_362_nl;
  wire and_1687_nl;
  wire and_1688_nl;
  wire mux_266_nl;
  wire mux_265_nl;
  wire mux_264_nl;
  wire or_391_nl;
  wire nor_246_nl;
  wire and_1697_nl;
  wire mux_551_nl;
  wire mux_550_nl;
  wire mux_549_nl;
  wire mux_548_nl;
  wire mux_547_nl;
  wire mux_546_nl;
  wire or_1135_nl;
  wire nor_486_nl;
  wire mux_545_nl;
  wire mux_544_nl;
  wire or_1136_nl;
  wire nor_487_nl;
  wire mux_543_nl;
  wire or_1137_nl;
  wire nor_488_nl;
  wire mux_542_nl;
  wire mux_541_nl;
  wire mux_540_nl;
  wire or_1138_nl;
  wire nor_489_nl;
  wire mux_539_nl;
  wire or_1139_nl;
  wire nor_490_nl;
  wire mux_538_nl;
  wire mux_537_nl;
  wire or_1140_nl;
  wire nor_491_nl;
  wire mux_536_nl;
  wire or_1141_nl;
  wire nor_492_nl;
  wire mux_535_nl;
  wire mux_534_nl;
  wire mux_533_nl;
  wire mux_532_nl;
  wire or_1142_nl;
  wire nor_493_nl;
  wire mux_531_nl;
  wire nand_47_nl;
  wire nor_494_nl;
  wire mux_530_nl;
  wire mux_529_nl;
  wire or_1143_nl;
  wire nor_495_nl;
  wire mux_528_nl;
  wire or_1144_nl;
  wire nor_496_nl;
  wire mux_527_nl;
  wire mux_526_nl;
  wire mux_525_nl;
  wire nand_48_nl;
  wire nor_497_nl;
  wire mux_524_nl;
  wire nand_49_nl;
  wire nor_498_nl;
  wire mux_523_nl;
  wire mux_522_nl;
  wire nand_50_nl;
  wire nor_499_nl;
  wire mux_521_nl;
  wire or_1145_nl;
  wire nor_500_nl;
  wire mux_520_nl;
  wire mux_519_nl;
  wire mux_518_nl;
  wire mux_517_nl;
  wire mux_516_nl;
  wire nand_51_nl;
  wire nor_501_nl;
  wire mux_515_nl;
  wire nand_52_nl;
  wire nor_502_nl;
  wire mux_514_nl;
  wire mux_513_nl;
  wire or_1146_nl;
  wire nor_503_nl;
  wire mux_512_nl;
  wire nand_53_nl;
  wire nor_504_nl;
  wire mux_511_nl;
  wire mux_510_nl;
  wire mux_509_nl;
  wire or_1147_nl;
  wire nor_505_nl;
  wire mux_508_nl;
  wire or_1148_nl;
  wire nor_506_nl;
  wire mux_507_nl;
  wire mux_506_nl;
  wire or_1149_nl;
  wire nor_507_nl;
  wire mux_505_nl;
  wire or_1150_nl;
  wire nor_508_nl;
  wire mux_504_nl;
  wire mux_503_nl;
  wire mux_502_nl;
  wire mux_501_nl;
  wire or_1151_nl;
  wire nor_509_nl;
  wire mux_500_nl;
  wire or_1152_nl;
  wire nor_510_nl;
  wire mux_499_nl;
  wire mux_498_nl;
  wire or_1153_nl;
  wire nor_511_nl;
  wire mux_497_nl;
  wire or_1154_nl;
  wire nor_512_nl;
  wire mux_496_nl;
  wire mux_495_nl;
  wire mux_494_nl;
  wire or_1155_nl;
  wire nor_513_nl;
  wire mux_493_nl;
  wire or_1156_nl;
  wire nor_514_nl;
  wire mux_492_nl;
  wire mux_491_nl;
  wire or_1157_nl;
  wire nor_515_nl;
  wire mux_490_nl;
  wire nand_54_nl;
  wire nor_516_nl;
  wire[6:0] MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[6:0] MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire[7:0] nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl;
  wire mux_724_nl;
  wire or_1188_nl;
  wire or_1191_nl;
  wire or_1192_nl;
  wire or_1193_nl;
  wire or_1194_nl;
  wire or_1195_nl;
  wire or_1196_nl;
  wire or_1197_nl;
  wire or_1198_nl;
  wire or_1199_nl;
  wire or_1200_nl;
  wire or_1201_nl;
  wire or_1219_nl;
  wire mux_741_nl;
  wire or_1216_nl;
  wire or_1220_nl;
  wire or_1221_nl;
  wire or_1222_nl;
  wire or_1223_nl;
  wire or_1224_nl;
  wire or_1225_nl;
  wire or_1226_nl;
  wire or_1227_nl;
  wire or_1228_nl;
  wire mux_752_nl;
  wire or_1229_nl;
  wire or_1231_nl;
  wire mux_759_nl;
  wire or_1246_nl;
  wire or_1251_nl;
  wire or_1252_nl;
  wire or_1253_nl;
  wire or_1254_nl;
  wire or_1255_nl;
  wire or_1256_nl;
  wire or_1257_nl;
  wire or_1258_nl;
  wire or_1259_nl;
  wire or_1260_nl;
  wire or_1262_nl;
  wire or_1261_nl;
  wire or_1263_nl;
  wire mux_772_nl;
  wire or_1281_nl;
  wire mux_781_nl;
  wire or_1277_nl;
  wire or_1282_nl;
  wire or_1283_nl;
  wire or_1284_nl;
  wire or_1285_nl;
  wire or_1286_nl;
  wire or_1287_nl;
  wire or_1288_nl;
  wire or_1289_nl;
  wire or_1290_nl;
  wire mux_793_nl;
  wire mux_792_nl;
  wire or_1291_nl;
  wire or_1292_nl;
  wire mux_796_nl;
  wire mux_795_nl;
  wire mux_824_nl;
  wire or_1309_nl;
  wire mux_825_nl;
  wire or_1333_nl;
  wire or_1335_nl;
  wire or_1336_nl;
  wire or_1337_nl;
  wire or_1338_nl;
  wire mux_831_nl;
  wire or_1339_nl;
  wire or_1341_nl;
  wire or_1342_nl;
  wire or_1343_nl;
  wire mux_835_nl;
  wire or_1344_nl;
  wire or_1346_nl;
  wire or_1362_nl;
  wire or_1360_nl;
  wire or_1363_nl;
  wire or_1364_nl;
  wire or_1365_nl;
  wire or_1366_nl;
  wire or_1367_nl;
  wire or_1368_nl;
  wire or_1369_nl;
  wire or_1370_nl;
  wire or_1371_nl;
  wire or_1372_nl;
  wire or_1374_nl;
  wire or_1373_nl;
  wire or_1375_nl;
  wire mux_852_nl;
  wire mux_856_nl;
  wire or_1388_nl;
  wire or_1390_nl;
  wire or_1391_nl;
  wire or_1392_nl;
  wire or_1393_nl;
  wire or_1394_nl;
  wire or_1395_nl;
  wire or_1396_nl;
  wire or_1397_nl;
  wire or_1398_nl;
  wire mux_868_nl;
  wire mux_867_nl;
  wire or_1399_nl;
  wire or_1400_nl;
  wire mux_871_nl;
  wire mux_870_nl;
  wire mux_904_nl;
  wire or_1439_nl;
  wire or_1440_nl;
  wire or_1441_nl;
  wire or_1442_nl;
  wire mux_910_nl;
  wire or_1443_nl;
  wire or_1445_nl;
  wire or_1446_nl;
  wire or_1447_nl;
  wire mux_914_nl;
  wire or_1448_nl;
  wire or_1450_nl;
  wire or_1463_nl;
  wire or_1464_nl;
  wire or_1465_nl;
  wire or_1466_nl;
  wire or_1467_nl;
  wire or_1468_nl;
  wire or_1469_nl;
  wire or_1470_nl;
  wire or_1471_nl;
  wire or_1472_nl;
  wire or_1474_nl;
  wire or_1473_nl;
  wire or_1475_nl;
  wire mux_931_nl;
  wire or_1487_nl;
  wire or_1488_nl;
  wire or_1489_nl;
  wire or_1490_nl;
  wire or_1491_nl;
  wire or_1492_nl;
  wire or_1493_nl;
  wire or_1494_nl;
  wire or_1495_nl;
  wire mux_946_nl;
  wire mux_945_nl;
  wire or_1496_nl;
  wire or_1497_nl;
  wire mux_949_nl;
  wire mux_948_nl;
  wire or_1531_nl;
  wire mux_1112_nl;
  wire mux_1117_nl;
  wire or_1542_nl;
  wire or_1543_nl;
  wire or_1544_nl;
  wire or_1545_nl;
  wire mux_988_nl;
  wire or_1546_nl;
  wire or_1548_nl;
  wire or_1549_nl;
  wire or_1550_nl;
  wire mux_993_nl;
  wire mux_992_nl;
  wire or_1551_nl;
  wire mux_996_nl;
  wire mux_995_nl;
  wire mux_983_nl;
  wire mux_1113_nl;
  wire mux_1039_nl;
  wire mux_319_nl;
  wire mux_318_nl;
  wire or_242_nl;
  wire mux_395_nl;
  wire mux_394_nl;
  wire mux_393_nl;
  wire mux_392_nl;
  wire mux_391_nl;
  wire mux_390_nl;
  wire mux_389_nl;
  wire or_563_nl;
  wire or_562_nl;
  wire mux_388_nl;
  wire mux_387_nl;
  wire mux_386_nl;
  wire nor_371_nl;
  wire mux_385_nl;
  wire mux_384_nl;
  wire nor_373_nl;
  wire mux_383_nl;
  wire mux_382_nl;
  wire mux_381_nl;
  wire or_553_nl;
  wire or_552_nl;
  wire mux_380_nl;
  wire or_551_nl;
  wire or_550_nl;
  wire mux_379_nl;
  wire mux_378_nl;
  wire mux_377_nl;
  wire nor_375_nl;
  wire mux_376_nl;
  wire or_545_nl;
  wire or_544_nl;
  wire mux_375_nl;
  wire mux_374_nl;
  wire mux_373_nl;
  wire mux_372_nl;
  wire mux_371_nl;
  wire nor_377_nl;
  wire mux_370_nl;
  wire or_539_nl;
  wire or_538_nl;
  wire mux_369_nl;
  wire mux_368_nl;
  wire or_537_nl;
  wire or_536_nl;
  wire mux_367_nl;
  wire or_535_nl;
  wire or_534_nl;
  wire mux_366_nl;
  wire mux_365_nl;
  wire mux_364_nl;
  wire mux_363_nl;
  wire nor_379_nl;
  wire mux_362_nl;
  wire or_529_nl;
  wire or_528_nl;
  wire mux_361_nl;
  wire mux_360_nl;
  wire or_527_nl;
  wire or_526_nl;
  wire mux_359_nl;
  wire or_525_nl;
  wire or_524_nl;
  wire mux_358_nl;
  wire mux_357_nl;
  wire mux_356_nl;
  wire mux_355_nl;
  wire mux_354_nl;
  wire or_523_nl;
  wire or_522_nl;
  wire mux_353_nl;
  wire mux_352_nl;
  wire nor_381_nl;
  wire mux_351_nl;
  wire mux_350_nl;
  wire mux_349_nl;
  wire nor_383_nl;
  wire mux_348_nl;
  wire mux_347_nl;
  wire nor_385_nl;
  wire mux_346_nl;
  wire mux_345_nl;
  wire mux_344_nl;
  wire or_509_nl;
  wire or_508_nl;
  wire mux_343_nl;
  wire or_507_nl;
  wire or_506_nl;
  wire mux_342_nl;
  wire mux_341_nl;
  wire mux_340_nl;
  wire nor_387_nl;
  wire mux_339_nl;
  wire mux_338_nl;
  wire nor_389_nl;
  wire mux_337_nl;
  wire mux_336_nl;
  wire mux_335_nl;
  wire mux_334_nl;
  wire or_497_nl;
  wire or_496_nl;
  wire mux_333_nl;
  wire mux_332_nl;
  wire nor_391_nl;
  wire mux_331_nl;
  wire mux_330_nl;
  wire or_491_nl;
  wire or_490_nl;
  wire mux_329_nl;
  wire or_489_nl;
  wire and_578_nl;
  wire nor_70_nl;
  wire mux_328_nl;
  wire mux_327_nl;
  wire mux_326_nl;
  wire or_486_nl;
  wire or_485_nl;
  wire mux_325_nl;
  wire mux_324_nl;
  wire nor_393_nl;
  wire mux_323_nl;
  wire mux_322_nl;
  wire or_480_nl;
  wire or_479_nl;
  wire mux_321_nl;
  wire mux_320_nl;
  wire nor_394_nl;
  wire ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_64_nl;
  wire[4:0] and_1758_nl;
  wire[4:0] mux1h_1_nl;
  wire[4:0] MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[4:0] MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire[5:0] nl_MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl;
  wire and_1310_nl;
  wire or_1565_nl;
  wire mux_661_nl;
  wire nand_55_nl;
  wire or_1048_nl;
  wire mux_660_nl;
  wire mux_659_nl;
  wire mux_658_nl;
  wire or_1170_nl;
  wire nor_645_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_192_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_193_nl;
  wire and_1315_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_194_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_195_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_196_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_197_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_198_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_199_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_200_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_201_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_202_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_203_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_204_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_205_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_206_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_207_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_208_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_209_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_210_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_211_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_212_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_213_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_214_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_215_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_216_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_217_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_218_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_219_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_220_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_221_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_222_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_223_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_224_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_225_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_226_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_227_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_228_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_229_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_230_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_231_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_232_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_233_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_234_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_235_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_236_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_237_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_238_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_239_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_240_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_241_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_242_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_243_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_244_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_245_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_246_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_247_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_248_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_249_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_250_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_251_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_252_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_253_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_254_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_255_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_256_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_257_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_258_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_259_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_260_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_261_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_262_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_263_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_264_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_265_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_266_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_267_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_268_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_269_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_270_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_271_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_272_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_273_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_274_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_275_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_276_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_277_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_278_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_279_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_280_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_281_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_282_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_283_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_284_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_285_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_286_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_287_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_288_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_289_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_290_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_291_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_292_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_293_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_294_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_295_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_296_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_297_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_298_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_299_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_300_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_301_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_302_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_303_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_304_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_305_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_306_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_307_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_308_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_309_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_310_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_311_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_312_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_313_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_314_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_315_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_316_nl;
  wire result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_317_nl;
  wire not_2129_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl;
  wire[6:0] MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl;
  wire[6:0] MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire[7:0] nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl;
  wire and_1757_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_256_nl;
  wire[3:0] MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire[4:0] nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl;
  wire and_272_nl;
  wire result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_11_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_33_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl;
  wire[7:0] acc_nl;
  wire[8:0] nl_acc_nl;
  wire[6:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl;
  wire[4:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl;
  wire and_1939_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_322_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_323_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_98_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_318_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_319_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_99_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_320_nl;
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_321_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [12:0] nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , 1'b0};
  wire [12:0] nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl;
  wire [4:0] nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[4]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl
      = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      (MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg[3:0]), MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_1_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl;
  wire [5:0] nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl
      = MUX_v_4_2_2(MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1,
      (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva);
  assign nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_1_nl
      , MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_4_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_99_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_100_nl;
  wire [4:0] nl_MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_99_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg[4]), MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_100_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg[3:0]), MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_99_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_100_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_102_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_103_nl;
  wire [4:0] nl_MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_102_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg[4]), MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_103_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg[3:0]), MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_102_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_103_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_105_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_106_nl;
  wire [4:0] nl_MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_105_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[4]), MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_106_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg[3:0]), MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_105_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_106_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_108_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_109_nl;
  wire [4:0] nl_MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_108_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[4]), MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_109_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg[3:0]), MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_108_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_109_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_111_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_112_nl;
  wire [4:0] nl_MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_111_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg[4]), MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_112_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg[3:0]), MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_111_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_112_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_114_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_115_nl;
  wire [4:0] nl_MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_114_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg[4]), MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_115_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg[3:0]), MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_114_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_115_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_117_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_118_nl;
  wire [4:0] nl_MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_117_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg[4]), MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_118_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg[3:0]), MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_117_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_118_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_120_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_121_nl;
  wire [4:0] nl_MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_120_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg[4]), MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_121_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg[3:0]), MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_120_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_121_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_123_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_124_nl;
  wire [4:0] nl_MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_123_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[4]), MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_124_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg[3:0]), MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_123_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_124_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_126_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_127_nl;
  wire [4:0] nl_MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_126_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg[4]), MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_127_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg[3:0]), MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_126_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_127_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_129_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_130_nl;
  wire [4:0] nl_MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_129_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[4]), MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_130_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg[3:0]), MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_129_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_130_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_132_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_133_nl;
  wire [4:0] nl_MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_132_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg[4]), MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_133_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg[3:0]), MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_132_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_133_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_135_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_136_nl;
  wire [4:0] nl_MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_135_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[4]), MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_136_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg[3:0]), MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_135_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_136_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_138_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_139_nl;
  wire [4:0] nl_MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_138_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[4]), MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_139_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg[3:0]), MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_138_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_139_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_141_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_142_nl;
  wire [4:0] nl_MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_141_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[4]), MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_142_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg[3:0]), MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_141_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_142_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_144_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_145_nl;
  wire [4:0] nl_MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_144_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg[4]), MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_145_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg[3:0]), MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_144_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_145_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_147_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_148_nl;
  wire [4:0] nl_MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_147_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[4]), MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_148_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg[3:0]), MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_147_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_148_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_150_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_151_nl;
  wire [4:0] nl_MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_150_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[4]), MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_151_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg[3:0]), MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_150_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_151_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_153_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_154_nl;
  wire [4:0] nl_MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_153_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[4]), MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_154_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg[3:0]), MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_153_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_154_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_156_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_157_nl;
  wire [4:0] nl_MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_156_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg[4]), MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_157_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg[3:0]), MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_156_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_157_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_159_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_160_nl;
  wire [4:0] nl_MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_159_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[4]), MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_160_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg[3:0]), MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_159_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_160_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_162_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_163_nl;
  wire [4:0] nl_MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_162_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[4]), MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_163_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg[3:0]), MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_162_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_163_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_165_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_166_nl;
  wire [4:0] nl_MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_165_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[4]), MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_166_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg[3:0]), MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_165_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_166_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_168_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_169_nl;
  wire [4:0] nl_MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_168_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[4]), MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_169_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg[3:0]), MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_168_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_169_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_171_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_172_nl;
  wire [4:0] nl_MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_171_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[4]), MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_172_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg[3:0]), MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_171_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_172_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_174_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_175_nl;
  wire [4:0] nl_MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_174_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[4]), MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_175_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg[3:0]), MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_174_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_175_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_177_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_178_nl;
  wire [4:0] nl_MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_177_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[4]), MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_178_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg[3:0]), MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_177_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_178_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_180_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_181_nl;
  wire [4:0] nl_MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_180_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[4]), MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_181_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg[3:0]), MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_180_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_181_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_183_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_184_nl;
  wire [4:0] nl_MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_183_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[4]), MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_184_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg[3:0]), MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_183_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_184_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_186_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_187_nl;
  wire [4:0] nl_MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_186_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[4]), MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_187_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg[3:0]), MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_186_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_187_nl};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_189_nl;
  wire[3:0] ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_190_nl;
  wire [4:0] nl_MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_189_nl
      = MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[4]), MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_190_nl
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg[3:0]), MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign nl_MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_189_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_190_nl};
  wire [11:0] nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a;
  assign nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a = {operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 , 1'b0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl;
  wire [5:0] nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  assign nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_3_nl
      , MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl;
  wire [5:0] nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva;
  assign nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl;
  wire [5:0] nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva;
  assign nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_5_nl
      , MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl;
  wire [5:0] nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva;
  assign nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_6_nl
      , MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl;
  wire [5:0] nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva;
  assign nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_7_nl
      , MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl;
  wire [5:0] nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva;
  assign nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_8_nl
      , MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl;
  wire [5:0] nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  assign nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_9_nl
      , MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl;
  wire [5:0] nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  assign nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_10_nl
      , MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl;
  wire [5:0] nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  assign nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_11_nl
      , MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl;
  wire [5:0] nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva;
  assign nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_12_nl
      , MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl;
  wire [5:0] nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva;
  assign nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_13_nl
      , MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl;
  wire [5:0] nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva;
  assign nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_14_nl
      , MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl;
  wire [5:0] nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva;
  assign nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_15_nl
      , MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl;
  wire [5:0] nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva;
  assign nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_16_nl
      , MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_17_nl;
  wire [5:0] nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_17_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  assign nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_17_nl
      , MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_18_nl;
  wire [5:0] nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_18_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva;
  assign nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_18_nl
      , MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_19_nl;
  wire [5:0] nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_19_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva;
  assign nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_19_nl
      , MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_20_nl;
  wire [5:0] nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_20_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva;
  assign nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_20_nl
      , MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_21_nl;
  wire [5:0] nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_21_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva;
  assign nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_21_nl
      , MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_22_nl;
  wire [5:0] nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_22_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva;
  assign nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_22_nl
      , MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_23_nl;
  wire [5:0] nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_23_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva;
  assign nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_23_nl
      , MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_24_nl;
  wire [5:0] nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_24_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva;
  assign nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_24_nl
      , MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_25_nl;
  wire [5:0] nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_25_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva;
  assign nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_25_nl
      , MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_26_nl;
  wire [5:0] nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_26_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva;
  assign nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_26_nl
      , MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_27_nl;
  wire [5:0] nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_27_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva;
  assign nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_27_nl
      , MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_28_nl;
  wire [5:0] nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_28_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva;
  assign nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_28_nl
      , MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_29_nl;
  wire [5:0] nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_29_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva;
  assign nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_29_nl
      , MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_30_nl;
  wire [5:0] nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_30_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva;
  assign nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_30_nl
      , MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_31_nl;
  wire [5:0] nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_31_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva;
  assign nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_31_nl
      , MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_32_nl;
  wire [5:0] nl_MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_32_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1[0])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva;
  assign nl_MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_32_nl
      , MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm};
  wire [12:0] nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , 1'b0};
  wire ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl;
  wire [5:0] nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[1])
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva;
  assign nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s = {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_and_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm};
  wire [4:0] nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s;
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s
      = {1'b0, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva};
  wire [12:0] nl_MAC_52_leading_sign_13_1_1_0_rg_mantissa;
  assign nl_MAC_52_leading_sign_13_1_1_0_rg_mantissa = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  wire [12:0] nl_MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a;
  assign nl_MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a = {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 , (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])};
  ccs_in_v1 #(.rscid(32'sd1),
  .width(32'sd11)) input_m_rsci (
      .dat(input_m_rsc_dat),
      .idat(input_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd2),
  .width(32'sd5)) input_e_rsci (
      .dat(input_e_rsc_dat),
      .idat(input_e_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd3),
  .width(32'sd704)) taps_m_rsci (
      .dat(taps_m_rsc_dat),
      .idat(taps_m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd320)) taps_e_rsci (
      .dat(taps_e_rsc_dat),
      .idat(taps_e_rsci_idat)
    );
  ccs_out_v1 #(.rscid(32'sd5),
  .width(32'sd11)) return_m_rsci (
      .idat(return_m_rsci_idat),
      .dat(return_m_rsc_dat)
    );
  ccs_out_v1 #(.rscid(32'sd6),
  .width(32'sd5)) return_e_rsci (
      .idat(return_e_rsci_idat),
      .dat(return_e_rsc_dat)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_m_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(input_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) input_e_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(input_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_m_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(taps_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) taps_e_triosy_obj (
      .ld(reg_taps_e_triosy_obj_ld_cse),
      .lz(taps_e_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_m_triosy_obj (
      .ld(reg_return_e_triosy_obj_ld_cse),
      .lz(return_m_triosy_lz)
    );
  mgc_io_sync_v2 #(.valid(32'sd0)) return_e_triosy_obj (
      .ld(reg_return_e_triosy_obj_ld_cse),
      .lz(return_e_triosy_lz)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1),
      .z(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva),
      .s(nl_MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1),
      .z(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva),
      .s(nl_MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1),
      .z(MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva),
      .s(nl_MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1),
      .z(MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva),
      .s(nl_MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1),
      .z(MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva),
      .s(nl_MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1),
      .z(MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva),
      .s(nl_MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1),
      .z(MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva),
      .s(nl_MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1),
      .z(MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva),
      .s(nl_MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1),
      .z(MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva),
      .s(nl_MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1),
      .z(MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva),
      .s(nl_MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1),
      .z(MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva),
      .s(nl_MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1),
      .z(MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva),
      .s(nl_MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1),
      .z(MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva),
      .s(nl_MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1),
      .z(MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva),
      .s(nl_MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1),
      .z(MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva),
      .s(nl_MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1),
      .z(MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva),
      .s(nl_MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1),
      .z(MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva),
      .s(nl_MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1),
      .z(MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva),
      .s(nl_MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1),
      .z(MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva),
      .s(nl_MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1),
      .z(MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva),
      .s(nl_MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1),
      .z(MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva),
      .s(nl_MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1),
      .z(MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva),
      .s(nl_MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1),
      .z(MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva),
      .s(nl_MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1),
      .z(MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva),
      .s(nl_MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1),
      .z(MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva),
      .s(nl_MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1),
      .z(MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva),
      .s(nl_MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1),
      .z(MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva),
      .s(nl_MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1),
      .z(MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva),
      .s(nl_MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1),
      .z(MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva),
      .s(nl_MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1),
      .z(MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva),
      .s(nl_MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1),
      .z(MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva),
      .s(nl_MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1),
      .z(MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva),
      .s(nl_MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1),
      .z(MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva),
      .s(nl_MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[4:0]),
      .z(MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd12),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd12)) MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg (
      .a(nl_MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_rshift_rg_a[11:0]),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2),
      .z(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(nl_MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm),
      .z(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(nl_MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm),
      .z(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(nl_MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva),
      .s(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0),
      .z(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(nl_MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva),
      .s(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1),
      .z(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(nl_MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm),
      .z(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(nl_MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm),
      .z(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(nl_MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva),
      .z(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(nl_MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm),
      .z(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(nl_MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm),
      .z(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(nl_MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm),
      .z(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(nl_MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm),
      .z(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(nl_MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm),
      .z(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva),
      .s(nl_MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm),
      .z(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva),
      .s(nl_MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm),
      .z(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva),
      .s(nl_MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm),
      .z(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva),
      .s(nl_MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm),
      .z(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva),
      .s(nl_MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm),
      .z(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva),
      .s(nl_MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm),
      .z(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva),
      .s(nl_MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm),
      .z(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva),
      .s(nl_MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm),
      .z(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva),
      .s(nl_MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm),
      .z(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva),
      .s(nl_MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm),
      .z(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva),
      .s(nl_MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm),
      .z(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva),
      .s(nl_MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm),
      .z(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva),
      .s(nl_MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm),
      .z(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva),
      .s(nl_MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm),
      .z(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva),
      .s(nl_MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm),
      .z(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva),
      .s(nl_MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm),
      .z(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva),
      .s(nl_MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm),
      .z(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva),
      .s(nl_MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_r_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd4),
  .width_z(32'sd22)) MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva),
      .s(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm),
      .z(MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  leading_sign_13_1_1_0  MAC_1_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_1_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_54),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_56)
    );
  mgc_shift_l_v5 #(.width_a(32'sd22),
  .signd_a(32'sd0),
  .width_s(32'sd6),
  .width_z(32'sd22)) MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(nl_MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_rg_s[5:0]),
      .z(MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  mgc_shift_br_v5 #(.width_a(32'sd22),
  .signd_a(32'sd1),
  .width_s(32'sd5),
  .width_z(32'sd22)) MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg
      (
      .a(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva),
      .s(nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_rg_s[4:0]),
      .z(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm)
    );
  leading_sign_13_1_1_0  MAC_52_leading_sign_13_1_1_0_rg (
      .mantissa(nl_MAC_52_leading_sign_13_1_1_0_rg_mantissa[12:0]),
      .all_same(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_55),
      .rtn(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_57)
    );
  mgc_shift_l_v5 #(.width_a(32'sd13),
  .signd_a(32'sd0),
  .width_s(32'sd4),
  .width_z(32'sd13)) MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg (
      .a(nl_MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_rg_a[12:0]),
      .s(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0),
      .z(MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm)
    );
  fir_core_wait_dp fir_core_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg)
    );
  fir_core_core_fsm fir_core_core_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse = and_dcpl_105
      | and_dcpl_109;
  assign nor_459_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[4]));
  assign and_1670_cse = (fsm_output[4:3]==2'b11);
  assign nl_MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_39_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[199:195]);
  assign MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_91_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_116, and_1670_cse);
  assign or_1132_cse = (fsm_output[5]) | mux_91_nl;
  assign nor_457_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
      | (~ (fsm_output[1])));
  assign or_766_nl = (~ (fsm_output[0])) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6;
  assign mux_484_nl = MUX_s_1_2_2(nor_457_nl, (fsm_output[1]), or_766_nl);
  assign nor_458_nl = ~((fsm_output[6:2]!=5'b00000) | mux_484_nl);
  assign mux_485_nl = MUX_s_1_2_2(nor_458_nl, or_1132_cse, fsm_output[7]);
  assign or_770_rgt = mux_485_nl | (fsm_output[8]);
  assign and_930_rgt = (nor_459_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6)
      & and_dcpl_152 & and_dcpl_497;
  assign mux_159_nl = MUX_s_1_2_2(or_1120_cse, (~ or_1132_cse), fsm_output[7]);
  assign and_118_rgt = mux_159_nl & (~ (fsm_output[8]));
  assign nor_451_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[4]));
  assign or_224_cse = (fsm_output[3]) | (fsm_output[2]) | (fsm_output[1]) | (fsm_output[6]);
  assign nl_MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_38_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[194:190]);
  assign MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_85_nl = MUX_s_1_2_2((fsm_output[6]), or_224_cse, fsm_output[4]);
  assign or_1128_cse = (fsm_output[5]) | mux_85_nl;
  assign nor_449_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
      | (~ (fsm_output[1])));
  assign or_752_nl = (~ (fsm_output[0])) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6;
  assign mux_478_nl = MUX_s_1_2_2(nor_449_nl, (fsm_output[1]), or_752_nl);
  assign nor_450_nl = ~((fsm_output[6:2]!=5'b00000) | mux_478_nl);
  assign mux_479_nl = MUX_s_1_2_2(nor_450_nl, or_1128_cse, fsm_output[7]);
  assign or_756_rgt = mux_479_nl | (fsm_output[8]);
  assign and_922_rgt = (nor_451_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6)
      & and_dcpl_152 & and_dcpl_497;
  assign mux_161_nl = MUX_s_1_2_2(or_1120_cse, (~ or_1128_cse), fsm_output[7]);
  assign and_119_rgt = mux_161_nl & (~ (fsm_output[8]));
  assign and_1669_cse = (fsm_output[3:1]==3'b111);
  assign nor_447_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5);
  assign nl_MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_37_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[189:185]);
  assign MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_747_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[4]);
  assign mux_472_nl = MUX_s_1_2_2(nor_tmp_76, mux_tmp_468, or_747_nl);
  assign nor_77_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
      | (~ (fsm_output[0])));
  assign mux_473_nl = MUX_s_1_2_2(nor_tmp_76, mux_472_nl, nor_77_nl);
  assign mux_474_nl = MUX_s_1_2_2(mux_tmp_468, mux_473_nl, fsm_output[1]);
  assign mux_475_nl = MUX_s_1_2_2(mux_474_nl, nor_tmp_76, fsm_output[3]);
  assign and_1702_nl = (((fsm_output[3]) & (fsm_output[1])) | (fsm_output[6:4]!=3'b000))
      & (fsm_output[7]);
  assign mux_476_nl = MUX_s_1_2_2(mux_475_nl, and_1702_nl, fsm_output[2]);
  assign or_749_rgt = mux_476_nl | (fsm_output[8]);
  assign and_918_rgt = and_dcpl_152 & and_dcpl_259 & and_dcpl_85 & (nor_447_cse |
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6);
  assign nor_846_nl = ~((fsm_output[5:4]!=2'b00) | mux_tmp_159);
  assign mux_163_nl = MUX_s_1_2_2(or_1120_cse, nor_846_nl, fsm_output[7]);
  assign and_120_rgt = mux_163_nl & (~ (fsm_output[8]));
  assign nor_442_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5);
  assign or_741_cse = nor_442_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6;
  assign nl_MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_36_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[184:180]);
  assign MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_80_cse = MUX_s_1_2_2((fsm_output[6]), or_tmp_116, fsm_output[3]);
  assign or_1124_cse = (fsm_output[5:4]!=2'b00) | mux_80_cse;
  assign mux_468_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_741_cse);
  assign nor_443_nl = ~((fsm_output[5:2]!=4'b0000) | mux_468_nl);
  assign mux_469_nl = MUX_s_1_2_2(nor_443_nl, or_1124_cse, fsm_output[7]);
  assign or_743_rgt = mux_469_nl | (fsm_output[8]);
  assign and_913_rgt = and_dcpl_152 & or_741_cse & and_dcpl_497;
  assign mux_165_nl = MUX_s_1_2_2(or_1120_cse, (~ or_1124_cse), fsm_output[7]);
  assign and_121_rgt = mux_165_nl & (~ (fsm_output[8]));
  assign nor_438_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5);
  assign or_735_cse = nor_438_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6;
  assign nl_MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_35_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[179:175]);
  assign MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_465_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_735_cse);
  assign nor_439_nl = ~((fsm_output[5:2]!=4'b0000) | mux_465_nl);
  assign mux_466_nl = MUX_s_1_2_2(nor_439_nl, or_tmp_204, fsm_output[7]);
  assign or_737_rgt = mux_466_nl | (fsm_output[8]);
  assign and_909_rgt = and_dcpl_152 & or_735_cse & and_dcpl_497;
  assign mux_167_nl = MUX_s_1_2_2(or_1120_cse, (~ or_tmp_204), fsm_output[7]);
  assign and_122_rgt = mux_167_nl & (~ (fsm_output[8]));
  assign nor_434_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp[5:4]!=2'b00));
  assign or_1120_cse = (fsm_output[6:1]!=6'b000000);
  assign nl_MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_34_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[174:170]);
  assign MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nor_73_nl = ~(nor_434_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm));
  assign mux_462_nl = MUX_s_1_2_2(or_tmp_49, or_tmp_285, nor_73_nl);
  assign nor_435_nl = ~((fsm_output[5:2]!=4'b0000) | mux_462_nl);
  assign mux_463_nl = MUX_s_1_2_2(nor_435_nl, or_1120_cse, fsm_output[7]);
  assign or_729_rgt = mux_463_nl | (fsm_output[8]);
  assign and_905_rgt = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp[6])
      | nor_434_cse) & and_dcpl_152 & and_dcpl_497;
  assign nor_248_rgt = ~((~(or_1120_cse ^ (fsm_output[7]))) | (fsm_output[8]));
  assign nor_431_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp[5:4]!=2'b00));
  assign nl_MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_33_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[169:165]);
  assign MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nor_72_nl = ~(nor_431_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm));
  assign mux_459_nl = MUX_s_1_2_2(or_tmp_49, or_tmp_285, nor_72_nl);
  assign nor_432_nl = ~((fsm_output[4:2]!=3'b000) | mux_459_nl);
  assign mux_460_nl = MUX_s_1_2_2(nor_432_nl, nor_tmp_47, fsm_output[5]);
  assign or_723_rgt = mux_460_nl | or_dcpl_172;
  assign and_901_rgt = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp[6])
      | nor_431_cse) & and_dcpl_152 & and_dcpl_497;
  assign mux_168_nl = MUX_s_1_2_2(or_tmp_205, (~ nor_tmp_47), fsm_output[5]);
  assign and_125_rgt = mux_168_nl & and_dcpl_10;
  assign nor_428_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp[5:4]!=2'b00));
  assign nl_MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_32_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[164:160]);
  assign MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_715_nl = nor_428_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp[6]);
  assign mux_455_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_715_nl);
  assign mux_456_nl = MUX_s_1_2_2(or_tmp_49, mux_455_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm);
  assign nor_429_nl = ~((fsm_output[4:2]!=3'b000) | mux_456_nl);
  assign mux_457_nl = MUX_s_1_2_2(nor_429_nl, and_tmp_8, fsm_output[5]);
  assign or_717_rgt = mux_457_nl | or_dcpl_172;
  assign and_897_rgt = (nor_428_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_170_nl = MUX_s_1_2_2(or_tmp_205, (~ and_tmp_8), fsm_output[5]);
  assign and_127_rgt = mux_170_nl & and_dcpl_10;
  assign nor_425_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp[5:4]!=2'b00));
  assign nl_MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_31_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[159:155]);
  assign MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nor_71_nl = ~(nor_425_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm));
  assign mux_452_nl = MUX_s_1_2_2(or_tmp_49, or_tmp_285, nor_71_nl);
  assign nor_426_nl = ~((fsm_output[4:2]!=3'b000) | mux_452_nl);
  assign mux_453_nl = MUX_s_1_2_2(nor_426_nl, and_tmp_9, fsm_output[5]);
  assign or_710_rgt = mux_453_nl | or_dcpl_172;
  assign and_893_rgt = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp[6])
      | nor_425_cse) & and_dcpl_152 & and_dcpl_497;
  assign mux_172_nl = MUX_s_1_2_2(or_tmp_205, (~ and_tmp_9), fsm_output[5]);
  assign and_129_rgt = mux_172_nl & and_dcpl_10;
  assign nor_225_cse = ~((fsm_output[5]) | (fsm_output[7]));
  assign nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_30_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[154:150]);
  assign MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_450_nl = MUX_s_1_2_2((~ or_1164_cse), or_1164_cse, fsm_output[3]);
  assign or_703_nl = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[6])
      | (fsm_output[1:0]!=2'b01);
  assign mux_448_nl = MUX_s_1_2_2((fsm_output[1]), or_703_nl, fsm_output[2]);
  assign mux_449_nl = MUX_s_1_2_2((~ mux_448_nl), or_1164_cse, fsm_output[3]);
  assign or_702_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[5:4]!=2'b00);
  assign mux_451_nl = MUX_s_1_2_2(mux_450_nl, mux_449_nl, or_702_nl);
  assign or_704_rgt = mux_451_nl | or_dcpl_278;
  assign and_890_rgt = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp[5:4]!=2'b00))))
      & and_dcpl_158 & and_dcpl_547;
  assign and_133_rgt = (~((~(or_1164_cse ^ (fsm_output[3]))) | (fsm_output[8])))
      & and_dcpl_121;
  assign nor_421_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp[5:4]!=2'b00));
  assign nl_MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_29_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[149:145]);
  assign MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_695_nl = nor_421_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp[6]);
  assign mux_442_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_695_nl);
  assign mux_443_nl = MUX_s_1_2_2(or_tmp_49, mux_442_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm);
  assign nor_422_nl = ~((fsm_output[4:2]!=3'b000) | mux_443_nl);
  assign mux_444_nl = MUX_s_1_2_2(nor_422_nl, and_tmp_10, fsm_output[5]);
  assign or_697_rgt = mux_444_nl | or_dcpl_172;
  assign and_884_rgt = (nor_421_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_174_nl = MUX_s_1_2_2(or_tmp_205, (~ and_tmp_10), fsm_output[5]);
  assign and_135_rgt = mux_174_nl & and_dcpl_10;
  assign nor_415_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp[5:4]!=2'b00));
  assign nl_MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_28_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[144:140]);
  assign MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_680_nl = nor_415_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp[6]);
  assign mux_434_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_680_nl);
  assign or_681_nl = (fsm_output[3:2]!=2'b00) | mux_434_nl;
  assign mux_435_nl = MUX_s_1_2_2(or_224_cse, or_681_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm);
  assign nor_416_nl = ~((fsm_output[4]) | mux_435_nl);
  assign mux_436_nl = MUX_s_1_2_2(nor_416_nl, mux_tmp_172, fsm_output[5]);
  assign or_683_rgt = mux_436_nl | or_dcpl_172;
  assign and_876_rgt = (nor_415_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_176_nl = MUX_s_1_2_2(or_tmp_205, (~ mux_tmp_172), fsm_output[5]);
  assign and_137_rgt = mux_176_nl & and_dcpl_10;
  assign nor_412_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp[5:4]!=2'b00));
  assign nl_MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_27_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[139:135]);
  assign MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_177_nl = (fsm_output[4:3]!=2'b00);
  assign mux_59_cse = MUX_s_1_2_2(nor_tmp_7, (fsm_output[6]), or_177_nl);
  assign or_673_nl = nor_412_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp[6]);
  assign mux_430_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_673_nl);
  assign mux_431_nl = MUX_s_1_2_2(or_tmp_49, mux_430_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm);
  assign nor_413_nl = ~((fsm_output[4:2]!=3'b000) | mux_431_nl);
  assign mux_432_nl = MUX_s_1_2_2(nor_413_nl, mux_59_cse, fsm_output[5]);
  assign or_675_rgt = mux_432_nl | or_dcpl_172;
  assign and_872_rgt = (nor_412_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_178_nl = MUX_s_1_2_2(or_tmp_205, (~ mux_59_cse), fsm_output[5]);
  assign and_138_rgt = mux_178_nl & and_dcpl_10;
  assign nor_409_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp[5:4]!=2'b00));
  assign or_1113_cse = (fsm_output[4:1]!=4'b0000);
  assign nl_MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_26_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[134:130]);
  assign MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_665_nl = nor_409_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp[6]);
  assign mux_426_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_665_nl);
  assign mux_427_nl = MUX_s_1_2_2(or_tmp_49, mux_426_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm);
  assign nor_410_nl = ~((fsm_output[4:2]!=3'b000) | mux_427_nl);
  assign mux_428_nl = MUX_s_1_2_2(nor_410_nl, mux_tmp_176, fsm_output[5]);
  assign or_667_rgt = mux_428_nl | or_dcpl_172;
  assign and_868_rgt = (nor_409_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_180_nl = MUX_s_1_2_2(or_tmp_205, (~ mux_tmp_176), fsm_output[5]);
  assign and_139_rgt = mux_180_nl & and_dcpl_10;
  assign nor_406_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp[5:4]!=2'b00));
  assign nl_MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_25_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[129:125]);
  assign MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_657_nl = nor_406_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp[6]);
  assign mux_420_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_657_nl);
  assign or_658_nl = (fsm_output[2]) | mux_420_nl;
  assign mux_421_nl = MUX_s_1_2_2(or_tmp_116, or_658_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm);
  assign nor_407_nl = ~((fsm_output[3]) | mux_421_nl);
  assign mux_422_nl = MUX_s_1_2_2(nor_407_nl, nor_tmp_10, fsm_output[4]);
  assign mux_423_nl = MUX_s_1_2_2(mux_422_nl, (fsm_output[6]), fsm_output[5]);
  assign or_660_rgt = mux_423_nl | or_dcpl_172;
  assign and_864_rgt = (nor_406_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_181_nl = MUX_s_1_2_2((~ or_224_cse), nor_tmp_10, fsm_output[4]);
  assign mux_182_nl = MUX_s_1_2_2(mux_181_nl, (fsm_output[6]), fsm_output[5]);
  assign and_140_rgt = (~ mux_182_nl) & and_dcpl_10;
  assign nor_403_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp[5:4]!=2'b00));
  assign nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_24_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[124:120]);
  assign MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_651_nl = nor_403_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp[6]);
  assign mux_414_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_651_nl);
  assign mux_415_nl = MUX_s_1_2_2(or_tmp_49, mux_414_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm);
  assign nor_404_nl = ~((fsm_output[3:2]!=2'b00) | mux_415_nl);
  assign mux_416_nl = MUX_s_1_2_2(nor_404_nl, and_tmp_11, fsm_output[4]);
  assign mux_417_nl = MUX_s_1_2_2(mux_416_nl, (fsm_output[6]), fsm_output[5]);
  assign or_653_rgt = mux_417_nl | or_dcpl_172;
  assign and_860_rgt = (nor_403_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_183_nl = MUX_s_1_2_2((~ or_224_cse), and_tmp_11, fsm_output[4]);
  assign mux_184_nl = MUX_s_1_2_2(mux_183_nl, (fsm_output[6]), fsm_output[5]);
  assign and_141_rgt = (~ mux_184_nl) & and_dcpl_10;
  assign nor_401_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp[5:4]!=2'b00));
  assign nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_23_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[119:115]);
  assign MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_644_nl = nor_401_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp[6]);
  assign mux_408_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_644_nl);
  assign or_645_nl = (fsm_output[3:2]!=2'b00) | mux_408_nl;
  assign mux_409_nl = MUX_s_1_2_2(or_224_cse, or_645_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm);
  assign mux_410_nl = MUX_s_1_2_2((~ mux_409_nl), mux_tmp_44, fsm_output[4]);
  assign mux_411_nl = MUX_s_1_2_2(mux_410_nl, (fsm_output[6]), fsm_output[5]);
  assign or_646_rgt = mux_411_nl | or_dcpl_172;
  assign and_856_rgt = (nor_401_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_185_nl = MUX_s_1_2_2((~ or_224_cse), mux_tmp_44, fsm_output[4]);
  assign mux_186_nl = MUX_s_1_2_2(mux_185_nl, (fsm_output[6]), fsm_output[5]);
  assign and_142_rgt = (~ mux_186_nl) & and_dcpl_10;
  assign nor_398_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp[5:4]!=2'b00));
  assign nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_22_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[114:110]);
  assign MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_637_nl = nor_398_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp[6]);
  assign mux_402_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_637_nl);
  assign mux_403_nl = MUX_s_1_2_2(or_tmp_49, mux_402_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm);
  assign nor_399_nl = ~((fsm_output[3:2]!=2'b00) | mux_403_nl);
  assign mux_404_nl = MUX_s_1_2_2(nor_399_nl, mux_tmp_170, fsm_output[4]);
  assign mux_405_nl = MUX_s_1_2_2(mux_404_nl, (fsm_output[6]), fsm_output[5]);
  assign or_639_rgt = mux_405_nl | or_dcpl_172;
  assign and_852_rgt = (nor_398_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_187_nl = MUX_s_1_2_2((~ or_224_cse), mux_tmp_170, fsm_output[4]);
  assign mux_188_nl = MUX_s_1_2_2(mux_187_nl, (fsm_output[6]), fsm_output[5]);
  assign and_143_rgt = (~ mux_188_nl) & and_dcpl_10;
  assign nor_396_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp[5:4]!=2'b00));
  assign or_627_cse = (fsm_output[5:4]!=2'b00);
  assign nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_21_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[109:105]);
  assign MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_629_nl = nor_396_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp[6]);
  assign mux_396_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_629_nl);
  assign or_630_nl = (fsm_output[2]) | mux_396_nl;
  assign mux_397_nl = MUX_s_1_2_2(or_tmp_116, or_630_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm);
  assign mux_398_nl = MUX_s_1_2_2((~ mux_397_nl), nor_tmp_7, fsm_output[3]);
  assign mux_399_nl = MUX_s_1_2_2(mux_398_nl, (fsm_output[6]), or_627_cse);
  assign or_631_rgt = mux_399_nl | or_dcpl_172;
  assign and_848_rgt = (nor_396_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_189_nl = MUX_s_1_2_2((~ or_tmp_116), nor_tmp_7, fsm_output[3]);
  assign mux_190_nl = MUX_s_1_2_2(mux_189_nl, (fsm_output[6]), or_627_cse);
  assign and_144_rgt = (~ mux_190_nl) & and_dcpl_10;
  assign nor_68_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign or_150_cse = (fsm_output[7]) | (fsm_output[5]) | (fsm_output[4]) | (fsm_output[3]);
  assign and_1698_cse = (fsm_output[1:0]==2'b11);
  assign or_151_cse = (~ (fsm_output[1])) | (fsm_output[0]) | (fsm_output[8]);
  assign or_152_cse = (fsm_output[6]) | (fsm_output[8]);
  assign nor_369_cse = ~((MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_20_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[104:100]);
  assign MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_192_nl = MUX_s_1_2_2(or_tmp_213, or_151_cse, fsm_output[6]);
  assign or_326_nl = and_1698_cse | (fsm_output[8]);
  assign mux_191_nl = MUX_s_1_2_2(or_326_nl, or_151_cse, fsm_output[6]);
  assign mux_193_nl = MUX_s_1_2_2(mux_192_nl, mux_191_nl, fsm_output[2]);
  assign mux_194_itm = MUX_s_1_2_2(mux_193_nl, or_151_cse, or_150_cse);
  assign nor_364_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp[5:4]!=2'b00));
  assign nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_19_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[99:95]);
  assign MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_468_nl = nor_364_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp[6]);
  assign mux_311_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_468_nl);
  assign mux_312_nl = MUX_s_1_2_2(or_tmp_49, mux_311_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm);
  assign nor_365_nl = ~((fsm_output[2]) | mux_312_nl);
  assign mux_313_nl = MUX_s_1_2_2(nor_365_nl, mux_tmp_166, fsm_output[3]);
  assign mux_314_nl = MUX_s_1_2_2(mux_313_nl, (fsm_output[6]), or_627_cse);
  assign or_470_rgt = mux_314_nl | or_dcpl_172;
  assign and_559_rgt = (nor_364_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_195_nl = MUX_s_1_2_2((~ or_tmp_116), mux_tmp_166, fsm_output[3]);
  assign mux_196_nl = MUX_s_1_2_2(mux_195_nl, (fsm_output[6]), or_627_cse);
  assign and_145_rgt = (~ mux_196_nl) & and_dcpl_10;
  assign or_452_cse = (fsm_output[4:2]!=3'b000);
  assign nor_360_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[5:4]!=2'b00));
  assign or_456_cse = (fsm_output[5:2]!=4'b0000);
  assign nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_18_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[94:90]);
  assign MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_301_nl = MUX_s_1_2_2(mux_tmp_294, (fsm_output[6]), or_452_cse);
  assign mux_298_nl = MUX_s_1_2_2(or_tmp_213, (fsm_output[1]), fsm_output[6]);
  assign or_451_nl = nor_360_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[6]);
  assign mux_299_nl = MUX_s_1_2_2(mux_298_nl, mux_tmp_294, or_451_nl);
  assign mux_300_nl = MUX_s_1_2_2(mux_299_nl, (fsm_output[6]), or_452_cse);
  assign mux_302_nl = MUX_s_1_2_2(mux_301_nl, mux_300_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_303_nl = MUX_s_1_2_2(mux_302_nl, (fsm_output[6]), fsm_output[5]);
  assign or_453_rgt = mux_303_nl | or_dcpl_172;
  assign and_551_rgt = (nor_360_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign and_146_rgt = ((or_dcpl_115 | or_627_cse) ^ (fsm_output[6])) & and_dcpl_10;
  assign nor_357_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[5:4]!=2'b00));
  assign nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_17_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[89:85]);
  assign MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_442_nl = nor_357_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[6]);
  assign mux_293_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_442_nl);
  assign or_443_nl = (fsm_output[2]) | mux_293_nl;
  assign mux_294_nl = MUX_s_1_2_2(or_1164_cse, or_443_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm);
  assign nor_358_nl = ~((fsm_output[4:3]!=2'b00) | mux_294_nl);
  assign mux_295_nl = MUX_s_1_2_2(nor_358_nl, nor_tmp_53, fsm_output[5]);
  assign or_445_rgt = mux_295_nl | or_dcpl_150;
  assign and_547_rgt = (nor_357_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_197_nl = MUX_s_1_2_2(or_1113_cse, (~ nor_tmp_53), fsm_output[5]);
  assign and_149_rgt = mux_197_nl & and_dcpl_2;
  assign nor_354_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[5:4]!=2'b00));
  assign nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_16_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[84:80]);
  assign MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_435_nl = nor_354_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[6]);
  assign mux_289_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_435_nl);
  assign mux_290_nl = MUX_s_1_2_2((fsm_output[1]), mux_289_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm);
  assign nor_355_nl = ~((fsm_output[4:2]!=3'b000) | mux_290_nl);
  assign mux_291_nl = MUX_s_1_2_2(nor_355_nl, and_tmp_12, fsm_output[5]);
  assign or_437_rgt = mux_291_nl | or_dcpl_150;
  assign and_543_rgt = (nor_354_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_198_nl = MUX_s_1_2_2(or_1113_cse, (~ and_tmp_12), fsm_output[5]);
  assign and_151_rgt = mux_198_nl & and_dcpl_2;
  assign nor_351_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[5:4]!=2'b00));
  assign nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_15_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[79:75]);
  assign MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_123_cse = (fsm_output[3]) | nor_tmp;
  assign and_1700_nl = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      & (fsm_output[0]))) & (fsm_output[1]);
  assign or_427_nl = nor_351_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[6]);
  assign mux_286_nl = MUX_s_1_2_2(and_1700_nl, (fsm_output[1]), or_427_nl);
  assign nor_352_nl = ~((fsm_output[4:2]!=3'b000) | mux_286_nl);
  assign mux_287_nl = MUX_s_1_2_2(nor_352_nl, and_tmp_13, fsm_output[5]);
  assign or_430_rgt = mux_287_nl | or_dcpl_150;
  assign and_539_rgt = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp[6])
      | nor_351_cse) & and_dcpl_152 & and_dcpl_497;
  assign mux_199_nl = MUX_s_1_2_2(or_1113_cse, (~ and_tmp_13), fsm_output[5]);
  assign and_153_rgt = mux_199_nl & and_dcpl_2;
  assign nor_348_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[5:4]!=2'b00));
  assign nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_14_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[74:70]);
  assign MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_420_nl = nor_348_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[6]);
  assign mux_282_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_420_nl);
  assign mux_283_nl = MUX_s_1_2_2((fsm_output[1]), mux_282_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign nor_349_nl = ~((fsm_output[4:2]!=3'b000) | mux_283_nl);
  assign mux_284_nl = MUX_s_1_2_2(nor_349_nl, and_tmp_14, fsm_output[5]);
  assign or_422_rgt = mux_284_nl | or_dcpl_150;
  assign and_535_rgt = (nor_348_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_200_nl = MUX_s_1_2_2(or_1113_cse, (~ and_tmp_14), fsm_output[5]);
  assign and_155_rgt = mux_200_nl & and_dcpl_2;
  assign nor_345_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[5:4]!=2'b00));
  assign nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_13_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[69:65]);
  assign MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_413_nl = nor_345_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[6]);
  assign mux_278_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_413_nl);
  assign mux_279_nl = MUX_s_1_2_2((fsm_output[1]), mux_278_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign nor_346_nl = ~((fsm_output[4:2]!=3'b000) | mux_279_nl);
  assign mux_280_nl = MUX_s_1_2_2(nor_346_nl, or_tmp_217, fsm_output[5]);
  assign or_415_rgt = mux_280_nl | or_dcpl_150;
  assign and_531_rgt = (nor_345_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_201_nl = MUX_s_1_2_2(or_1113_cse, (~ or_tmp_217), fsm_output[5]);
  assign and_156_rgt = mux_201_nl & and_dcpl_2;
  assign nor_342_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[5:4]!=2'b00));
  assign nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_12_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[64:60]);
  assign MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign and_4_cse = (fsm_output[3]) & or_1164_cse;
  assign or_406_nl = nor_342_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[6]);
  assign mux_274_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_406_nl);
  assign mux_275_nl = MUX_s_1_2_2((fsm_output[1]), mux_274_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign nor_343_nl = ~((fsm_output[4:2]!=3'b000) | mux_275_nl);
  assign mux_276_nl = MUX_s_1_2_2(nor_343_nl, or_tmp_218, fsm_output[5]);
  assign or_408_rgt = mux_276_nl | or_dcpl_150;
  assign and_527_rgt = (nor_342_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_202_nl = MUX_s_1_2_2(or_1113_cse, (~ or_tmp_218), fsm_output[5]);
  assign and_158_rgt = mux_202_nl & and_dcpl_2;
  assign nor_339_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[5:4]!=2'b00));
  assign nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_11_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[59:55]);
  assign MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_399_nl = nor_339_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[6]);
  assign mux_270_nl = MUX_s_1_2_2((~ or_tmp_213), (fsm_output[1]), or_399_nl);
  assign mux_271_nl = MUX_s_1_2_2((fsm_output[1]), mux_270_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm);
  assign nor_340_nl = ~((fsm_output[4:2]!=3'b000) | mux_271_nl);
  assign mux_272_nl = MUX_s_1_2_2(nor_340_nl, or_tmp_6, fsm_output[5]);
  assign or_401_rgt = mux_272_nl | or_dcpl_150;
  assign and_523_rgt = (nor_339_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_203_nl = MUX_s_1_2_2(or_1113_cse, (~ or_tmp_6), fsm_output[5]);
  assign and_159_rgt = mux_203_nl & and_dcpl_2;
  assign nor_455_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[4]));
  assign nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_1_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[14:10]);
  assign MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign nor_453_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
      | (~ (fsm_output[1])));
  assign or_759_nl = (~ (fsm_output[0])) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6;
  assign mux_481_nl = MUX_s_1_2_2(nor_453_nl, (fsm_output[1]), or_759_nl);
  assign nor_454_nl = ~((fsm_output[6:2]!=5'b00000) | mux_481_nl);
  assign mux_482_nl = MUX_s_1_2_2(nor_454_nl, or_tmp_222, fsm_output[7]);
  assign or_763_rgt = mux_482_nl | (fsm_output[8]);
  assign and_926_rgt = (nor_455_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6)
      & and_dcpl_152 & and_dcpl_497;
  assign mux_205_nl = MUX_s_1_2_2(or_1120_cse, (~ or_tmp_222), fsm_output[7]);
  assign and_160_rgt = mux_205_nl & (~ (fsm_output[8]));
  assign nor_418_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp[5:4]!=2'b00));
  assign nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(delay_lane_e_0_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[9:5]);
  assign MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign mux_65_cse = MUX_s_1_2_2(nor_tmp_10, (fsm_output[6]), fsm_output[4]);
  assign or_688_nl = nor_418_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp[6]);
  assign mux_438_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_688_nl);
  assign mux_439_nl = MUX_s_1_2_2(or_tmp_49, mux_438_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm);
  assign nor_419_nl = ~((fsm_output[4:2]!=3'b000) | mux_439_nl);
  assign mux_440_nl = MUX_s_1_2_2(nor_419_nl, mux_65_cse, fsm_output[5]);
  assign or_690_rgt = mux_440_nl | or_dcpl_172;
  assign and_880_rgt = (nor_418_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_207_nl = MUX_s_1_2_2(or_tmp_205, (~ mux_65_cse), fsm_output[5]);
  assign and_161_rgt = mux_207_nl & and_dcpl_10;
  assign nor_362_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp[5:4]!=2'b00));
  assign or_458_cse = (fsm_output[5:3]!=3'b000);
  assign nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = conv_s2s_5_6(input_e_rsci_idat)
      + conv_s2s_5_6(taps_e_rsci_idat[4:0]);
  assign MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm = nl_MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5:0];
  assign or_460_nl = nor_362_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp[6]);
  assign mux_305_nl = MUX_s_1_2_2(or_tmp_285, or_tmp_49, or_460_nl);
  assign mux_306_nl = MUX_s_1_2_2(or_tmp_49, mux_305_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_307_nl = MUX_s_1_2_2((~ mux_306_nl), nor_tmp_49, fsm_output[2]);
  assign mux_308_nl = MUX_s_1_2_2(mux_307_nl, (fsm_output[6]), or_458_cse);
  assign or_462_rgt = mux_308_nl | or_dcpl_172;
  assign and_555_rgt = (nor_362_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm))
      & and_dcpl_152 & and_dcpl_497;
  assign mux_208_nl = MUX_s_1_2_2((~ or_tmp_49), nor_tmp_49, fsm_output[2]);
  assign mux_209_nl = MUX_s_1_2_2(mux_208_nl, (fsm_output[6]), or_458_cse);
  assign and_162_rgt = (~ mux_209_nl) & and_dcpl_10;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
      = (~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_151;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse
      = MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_151;
  assign or_351_cse = (fsm_output[7:2]!=6'b000000);
  assign and_1312_m1c = and_dcpl_919 & and_dcpl_101;
  assign and_1317_m1c = and_dcpl_108 & and_dcpl_1287;
  assign and_1318_m1c = and_dcpl_919 & and_dcpl_1287;
  assign and_1321_m1c = and_dcpl_108 & and_dcpl_1291;
  assign and_1322_m1c = and_dcpl_919 & and_dcpl_1291;
  assign and_1325_m1c = and_dcpl_108 & and_dcpl_1295;
  assign and_1326_m1c = and_dcpl_919 & and_dcpl_1295;
  assign and_1328_m1c = and_dcpl_108 & and_dcpl_1298;
  assign and_1329_m1c = and_dcpl_919 & and_dcpl_1298;
  assign and_1331_m1c = and_dcpl_108 & and_dcpl_1301;
  assign and_1332_m1c = and_dcpl_919 & and_dcpl_1301;
  assign and_1334_m1c = and_dcpl_108 & and_dcpl_1304;
  assign and_1335_m1c = and_dcpl_919 & and_dcpl_1304;
  assign and_1337_m1c = and_dcpl_108 & and_dcpl_1307;
  assign and_1338_m1c = and_dcpl_919 & and_dcpl_1307;
  assign and_1339_m1c = and_dcpl_1006 & and_dcpl_101;
  assign and_1340_m1c = and_dcpl_1101 & and_dcpl_101;
  assign and_1341_m1c = and_dcpl_1006 & and_dcpl_1287;
  assign and_1342_m1c = and_dcpl_1101 & and_dcpl_1287;
  assign and_1343_m1c = and_dcpl_1006 & and_dcpl_1291;
  assign and_1344_m1c = and_dcpl_1101 & and_dcpl_1291;
  assign and_1345_m1c = and_dcpl_1006 & and_dcpl_1295;
  assign and_1346_m1c = and_dcpl_1101 & and_dcpl_1295;
  assign and_1347_m1c = and_dcpl_1006 & and_dcpl_1298;
  assign and_1348_m1c = and_dcpl_1101 & and_dcpl_1298;
  assign and_1349_m1c = and_dcpl_1006 & and_dcpl_1301;
  assign and_1350_m1c = and_dcpl_1101 & and_dcpl_1301;
  assign and_1351_m1c = and_dcpl_1006 & and_dcpl_1304;
  assign and_1352_m1c = and_dcpl_1101 & and_dcpl_1304;
  assign and_1353_m1c = and_dcpl_1006 & and_dcpl_1307;
  assign and_1354_m1c = and_dcpl_1101 & and_dcpl_1307;
  assign and_1356_m1c = and_dcpl_108 & and_dcpl_1326;
  assign and_1357_m1c = and_dcpl_919 & and_dcpl_1326;
  assign and_1359_m1c = and_dcpl_108 & and_dcpl_1329;
  assign and_1360_m1c = and_dcpl_919 & and_dcpl_1329;
  assign and_1362_m1c = and_dcpl_108 & and_dcpl_1332;
  assign and_1363_m1c = and_dcpl_919 & and_dcpl_1332;
  assign and_1365_m1c = and_dcpl_108 & and_dcpl_1335;
  assign and_1366_m1c = and_dcpl_919 & and_dcpl_1335;
  assign and_1368_m1c = and_dcpl_108 & and_dcpl_1338;
  assign and_1369_m1c = and_dcpl_919 & and_dcpl_1338;
  assign and_1371_m1c = and_dcpl_108 & and_dcpl_1341;
  assign and_1372_m1c = and_dcpl_919 & and_dcpl_1341;
  assign and_1374_m1c = and_dcpl_108 & and_dcpl_1344;
  assign and_1375_m1c = and_dcpl_919 & and_dcpl_1344;
  assign and_1377_m1c = and_dcpl_108 & and_dcpl_1347;
  assign and_1378_m1c = and_dcpl_919 & and_dcpl_1347;
  assign and_1379_m1c = and_dcpl_1006 & and_dcpl_1326;
  assign and_1380_m1c = and_dcpl_1101 & and_dcpl_1326;
  assign and_1381_m1c = and_dcpl_1006 & and_dcpl_1329;
  assign and_1382_m1c = and_dcpl_1101 & and_dcpl_1329;
  assign and_1383_m1c = and_dcpl_1006 & and_dcpl_1332;
  assign and_1384_m1c = and_dcpl_1101 & and_dcpl_1332;
  assign and_1385_m1c = and_dcpl_1006 & and_dcpl_1335;
  assign and_1386_m1c = and_dcpl_1101 & and_dcpl_1335;
  assign and_1387_m1c = and_dcpl_1006 & and_dcpl_1338;
  assign and_1388_m1c = and_dcpl_1101 & and_dcpl_1338;
  assign and_1389_m1c = and_dcpl_1006 & and_dcpl_1341;
  assign and_1390_m1c = and_dcpl_1101 & and_dcpl_1341;
  assign and_1391_m1c = and_dcpl_1006 & and_dcpl_1344;
  assign and_1392_m1c = and_dcpl_1101 & and_dcpl_1344;
  assign and_1393_m1c = and_dcpl_1006 & and_dcpl_1347;
  assign and_1394_m1c = and_dcpl_1101 & and_dcpl_1347;
  assign and_1829_cse = and_dcpl_1335 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm;
  assign mux_1035_itm = MUX_s_1_2_2(mux_tmp_976, or_tmp_746, and_1829_cse);
  assign and_1827_cse = and_dcpl_1335 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm;
  assign mux_1020_nl = MUX_s_1_2_2(mux_tmp_1010, mux_tmp_1009, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign mux_1021_nl = MUX_s_1_2_2(mux_tmp_994, mux_1020_nl, and_dcpl_1326);
  assign mux_1017_nl = MUX_s_1_2_2(mux_tmp_994, mux_1035_itm, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_1110_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_1016_nl = MUX_s_1_2_2(mux_1110_nl, or_tmp_746, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_1018_nl = MUX_s_1_2_2(mux_1017_nl, mux_1016_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_1014_nl = MUX_s_1_2_2(mux_tmp_1010, mux_tmp_1009, or_tmp_776);
  assign mux_1114_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_1011_nl = MUX_s_1_2_2(mux_1114_nl, or_tmp_746, or_tmp_776);
  assign mux_1015_nl = MUX_s_1_2_2(mux_1014_nl, mux_1011_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_1019_nl = MUX_s_1_2_2(mux_1018_nl, mux_1015_nl, and_dcpl_1326);
  assign mux_1022_nl = MUX_s_1_2_2(mux_1021_nl, mux_1019_nl, and_dcpl_1329);
  assign mux_1008_nl = MUX_s_1_2_2(mux_tmp_996, mux_tmp_978, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign mux_1009_nl = MUX_s_1_2_2(mux_tmp_1001, mux_1008_nl, and_dcpl_1326);
  assign mux_1111_nl = MUX_s_1_2_2(mux_tmp_976, or_tmp_746, and_1829_cse);
  assign mux_1003_nl = MUX_s_1_2_2(mux_1111_nl, or_tmp_746, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_1005_nl = MUX_s_1_2_2(mux_tmp_1001, mux_1003_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_1115_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_1002_nl = MUX_s_1_2_2(mux_1115_nl, or_tmp_746, or_tmp_838);
  assign mux_1006_nl = MUX_s_1_2_2(mux_1005_nl, mux_1002_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_1000_nl = MUX_s_1_2_2(mux_tmp_996, mux_tmp_978, or_tmp_776);
  assign mux_1116_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_978_nl = MUX_s_1_2_2(mux_1116_nl, or_tmp_746, or_tmp_719);
  assign mux_1001_nl = MUX_s_1_2_2(mux_1000_nl, mux_978_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_1007_nl = MUX_s_1_2_2(mux_1006_nl, mux_1001_nl, and_dcpl_1326);
  assign mux_1010_nl = MUX_s_1_2_2(mux_1009_nl, mux_1007_nl, and_dcpl_1329);
  assign mux_1023_nl = MUX_s_1_2_2(mux_1022_nl, mux_1010_nl, and_dcpl_1341);
  assign mux_973_nl = MUX_s_1_2_2(mux_tmp_963, mux_tmp_962, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1507_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | mux_973_nl;
  assign mux_974_nl = MUX_s_1_2_2(mux_tmp_947, or_1507_nl, and_dcpl_1326);
  assign mux_970_nl = MUX_s_1_2_2(mux_tmp_947, mux_tmp_929, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_969_nl = MUX_s_1_2_2(mux_tmp_914, or_tmp_971, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_971_nl = MUX_s_1_2_2(mux_970_nl, mux_969_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_967_nl = MUX_s_1_2_2(mux_tmp_963, mux_tmp_962, or_tmp_776);
  assign mux_964_nl = MUX_s_1_2_2(mux_tmp_914, or_tmp_971, or_tmp_776);
  assign mux_968_nl = MUX_s_1_2_2(mux_967_nl, mux_964_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1505_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | mux_968_nl;
  assign mux_972_nl = MUX_s_1_2_2(mux_971_nl, or_1505_nl, and_dcpl_1326);
  assign or_1506_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
      | mux_972_nl;
  assign mux_975_nl = MUX_s_1_2_2(mux_974_nl, or_1506_nl, and_dcpl_1329);
  assign mux_961_nl = MUX_s_1_2_2(mux_tmp_949, mux_tmp_930, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1501_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | mux_961_nl;
  assign mux_962_nl = MUX_s_1_2_2(mux_tmp_954, or_1501_nl, and_dcpl_1326);
  assign mux_956_nl = MUX_s_1_2_2(mux_tmp_929, or_tmp_971, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_958_nl = MUX_s_1_2_2(mux_tmp_954, mux_956_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_955_nl = MUX_s_1_2_2(mux_tmp_914, or_tmp_971, or_tmp_838);
  assign mux_959_nl = MUX_s_1_2_2(mux_958_nl, mux_955_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_953_nl = MUX_s_1_2_2(mux_tmp_949, mux_tmp_930, or_tmp_776);
  assign mux_918_nl = MUX_s_1_2_2(mux_tmp_914, or_tmp_971, or_tmp_719);
  assign mux_954_nl = MUX_s_1_2_2(mux_953_nl, mux_918_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1498_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | mux_954_nl;
  assign mux_960_nl = MUX_s_1_2_2(mux_959_nl, or_1498_nl, and_dcpl_1326);
  assign or_1500_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
      | mux_960_nl;
  assign mux_963_nl = MUX_s_1_2_2(mux_962_nl, or_1500_nl, and_dcpl_1329);
  assign or_1502_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm
      | mux_963_nl;
  assign mux_976_nl = MUX_s_1_2_2(mux_975_nl, or_1502_nl, and_dcpl_1341);
  assign mux_1024_nl = MUX_s_1_2_2(mux_1023_nl, mux_976_nl, and_dcpl_1006);
  assign and_1749_nl = and_dcpl_108 & (and_dcpl_1344 | and_dcpl_1338 | and_dcpl_1298
      | and_dcpl_1287 | and_dcpl_1307 | and_dcpl_1291 | and_dcpl_1304 | and_dcpl_1332
      | and_dcpl_1295 | and_dcpl_1301 | and_dcpl_1347);
  assign or_1413_nl = and_dcpl_1344 | and_dcpl_1338 | and_dcpl_1298 | and_dcpl_1287
      | and_dcpl_101 | and_dcpl_1307 | and_dcpl_1291 | and_dcpl_1304 | and_dcpl_1332
      | and_dcpl_1295 | and_dcpl_1301 | and_dcpl_1347;
  assign mux_901_nl = MUX_s_1_2_2(and_1749_nl, or_1413_nl, and_dcpl_919);
  assign or_nl = and_dcpl_1341 | and_dcpl_1329 | and_dcpl_1326 | and_dcpl_1335;
  assign mux_1037_nl = MUX_s_1_2_2(mux_901_nl, or_tmp_746, or_nl);
  assign or_1563_nl = mux_1037_nl | and_dcpl_1006;
  assign mux_1025_nl = MUX_s_1_2_2(mux_1024_nl, or_1563_nl, MAC_3_result_operator_result_operator_nor_tmp);
  assign mux_895_nl = MUX_s_1_2_2(mux_tmp_885, mux_tmp_884, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1410_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
      | mux_895_nl;
  assign mux_896_nl = MUX_s_1_2_2(mux_tmp_869, or_1410_nl, and_dcpl_1326);
  assign mux_892_nl = MUX_s_1_2_2(mux_tmp_869, mux_tmp_850, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_891_nl = MUX_s_1_2_2(mux_tmp_835, or_tmp_864, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_893_nl = MUX_s_1_2_2(mux_892_nl, mux_891_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_889_nl = MUX_s_1_2_2(mux_tmp_885, mux_tmp_884, or_tmp_776);
  assign mux_886_nl = MUX_s_1_2_2(mux_tmp_835, or_tmp_864, or_tmp_776);
  assign mux_890_nl = MUX_s_1_2_2(mux_889_nl, mux_886_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1408_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
      | mux_890_nl;
  assign mux_894_nl = MUX_s_1_2_2(mux_893_nl, or_1408_nl, and_dcpl_1326);
  assign or_1409_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm
      | mux_894_nl;
  assign mux_897_nl = MUX_s_1_2_2(mux_896_nl, or_1409_nl, and_dcpl_1329);
  assign mux_883_nl = MUX_s_1_2_2(mux_tmp_871, mux_tmp_851, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1404_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
      | mux_883_nl;
  assign mux_884_nl = MUX_s_1_2_2(mux_tmp_876, or_1404_nl, and_dcpl_1326);
  assign mux_878_nl = MUX_s_1_2_2(mux_tmp_850, or_tmp_864, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_880_nl = MUX_s_1_2_2(mux_tmp_876, mux_878_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_877_nl = MUX_s_1_2_2(mux_tmp_835, or_tmp_864, or_tmp_838);
  assign mux_881_nl = MUX_s_1_2_2(mux_880_nl, mux_877_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_875_nl = MUX_s_1_2_2(mux_tmp_871, mux_tmp_851, or_tmp_776);
  assign mux_839_nl = MUX_s_1_2_2(mux_tmp_835, or_tmp_864, or_tmp_719);
  assign mux_876_nl = MUX_s_1_2_2(mux_875_nl, mux_839_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1401_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
      | mux_876_nl;
  assign mux_882_nl = MUX_s_1_2_2(mux_881_nl, or_1401_nl, and_dcpl_1326);
  assign or_1403_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm
      | mux_882_nl;
  assign mux_885_nl = MUX_s_1_2_2(mux_884_nl, or_1403_nl, and_dcpl_1329);
  assign or_1405_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
      | mux_885_nl;
  assign mux_898_nl = MUX_s_1_2_2(mux_897_nl, or_1405_nl, and_dcpl_1341);
  assign mux_820_nl = MUX_s_1_2_2(mux_tmp_810, mux_tmp_809, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1306_nl = or_tmp_718 | mux_820_nl;
  assign mux_821_nl = MUX_s_1_2_2(mux_tmp_794, or_1306_nl, and_dcpl_1326);
  assign mux_817_nl = MUX_s_1_2_2(mux_tmp_794, mux_tmp_770, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_816_nl = MUX_s_1_2_2(mux_tmp_752, mux_tmp_733, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_818_nl = MUX_s_1_2_2(mux_817_nl, mux_816_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_814_nl = MUX_s_1_2_2(mux_tmp_810, mux_tmp_809, or_tmp_776);
  assign mux_811_nl = MUX_s_1_2_2(mux_tmp_752, mux_tmp_733, or_tmp_776);
  assign mux_815_nl = MUX_s_1_2_2(mux_814_nl, mux_811_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1303_nl = or_tmp_718 | mux_815_nl;
  assign mux_819_nl = MUX_s_1_2_2(mux_818_nl, or_1303_nl, and_dcpl_1326);
  assign or_1304_nl = or_tmp_717 | mux_819_nl;
  assign mux_822_nl = MUX_s_1_2_2(mux_821_nl, or_1304_nl, and_dcpl_1329);
  assign mux_808_nl = MUX_s_1_2_2(mux_tmp_796, mux_tmp_771, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_1297_nl = or_tmp_718 | mux_808_nl;
  assign mux_809_nl = MUX_s_1_2_2(mux_tmp_801, or_1297_nl, and_dcpl_1326);
  assign mux_803_nl = MUX_s_1_2_2(mux_tmp_770, mux_tmp_733, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_805_nl = MUX_s_1_2_2(mux_tmp_801, mux_803_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva);
  assign mux_802_nl = MUX_s_1_2_2(mux_tmp_752, mux_tmp_733, or_tmp_838);
  assign mux_806_nl = MUX_s_1_2_2(mux_805_nl, mux_802_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign mux_800_nl = MUX_s_1_2_2(mux_tmp_796, mux_tmp_771, or_tmp_776);
  assign mux_756_nl = MUX_s_1_2_2(mux_tmp_752, mux_tmp_733, or_tmp_719);
  assign mux_801_nl = MUX_s_1_2_2(mux_800_nl, mux_756_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_1293_nl = or_tmp_718 | mux_801_nl;
  assign mux_807_nl = MUX_s_1_2_2(mux_806_nl, or_1293_nl, and_dcpl_1326);
  assign or_1295_nl = or_tmp_717 | mux_807_nl;
  assign mux_810_nl = MUX_s_1_2_2(mux_809_nl, or_1295_nl, and_dcpl_1329);
  assign or_1298_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm
      | mux_810_nl;
  assign mux_823_nl = MUX_s_1_2_2(mux_822_nl, or_1298_nl, and_dcpl_1341);
  assign mux_1038_nl = MUX_s_1_2_2(mux_898_nl, mux_823_nl, and_dcpl_1006);
  assign or_1564_nl = mux_1038_nl | MAC_3_result_operator_result_operator_nor_tmp;
  assign mux_1026_tmp = MUX_s_1_2_2(mux_1025_nl, or_1564_nl, and_dcpl_1101);
  assign MAC_10_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      & MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_10_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2,
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm
      = conv_s2s_6_7({MAC_10_r_ac_float_else_and_nl , MAC_10_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6:0];
  assign operator_13_2_true_AC_TRN_AC_WRAP_or_ssc = and_dcpl_105 | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1
      | and_dcpl_162 | and_dcpl_157;
  assign and_1740_nl = (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign nor_646_nl = ~((~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1102_nl = (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_718_nl = MUX_s_1_2_2(nor_646_nl, or_1102_nl, MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_719_nl = MUX_s_1_2_2(and_1740_nl, mux_718_nl, fsm_output[2]);
  assign nor_647_nl = ~((~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1100_nl = (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_716_nl = MUX_s_1_2_2(nor_647_nl, or_1100_nl, MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_648_nl = ~((~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1098_nl = (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_715_nl = MUX_s_1_2_2(nor_648_nl, or_1098_nl, MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_717_nl = MUX_s_1_2_2(mux_716_nl, mux_715_nl, fsm_output[2]);
  assign mux_720_nl = MUX_s_1_2_2(mux_719_nl, mux_717_nl, fsm_output[3]);
  assign nor_649_nl = ~((~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1096_nl = (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_712_nl = MUX_s_1_2_2(nor_649_nl, or_1096_nl, MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_650_nl = ~((~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1094_nl = (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_711_nl = MUX_s_1_2_2(nor_650_nl, or_1094_nl, MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_713_nl = MUX_s_1_2_2(mux_712_nl, mux_711_nl, fsm_output[2]);
  assign nor_651_nl = ~((~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1092_nl = (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_709_nl = MUX_s_1_2_2(nor_651_nl, or_1092_nl, MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_652_nl = ~((~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1090_nl = (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_708_nl = MUX_s_1_2_2(nor_652_nl, or_1090_nl, MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_710_nl = MUX_s_1_2_2(mux_709_nl, mux_708_nl, fsm_output[2]);
  assign mux_714_nl = MUX_s_1_2_2(mux_713_nl, mux_710_nl, fsm_output[3]);
  assign mux_721_nl = MUX_s_1_2_2(mux_720_nl, mux_714_nl, fsm_output[4]);
  assign nor_653_nl = ~((~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1088_nl = (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_704_nl = MUX_s_1_2_2(nor_653_nl, or_1088_nl, MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_1741_nl = (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1087_nl = (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_703_nl = MUX_s_1_2_2(and_1741_nl, or_1087_nl, MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_705_nl = MUX_s_1_2_2(mux_704_nl, mux_703_nl, fsm_output[2]);
  assign nor_654_nl = ~((~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1085_nl = (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_701_nl = MUX_s_1_2_2(nor_654_nl, or_1085_nl, MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_655_nl = ~((~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1083_nl = (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_700_nl = MUX_s_1_2_2(nor_655_nl, or_1083_nl, MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_702_nl = MUX_s_1_2_2(mux_701_nl, mux_700_nl, fsm_output[2]);
  assign mux_706_nl = MUX_s_1_2_2(mux_705_nl, mux_702_nl, fsm_output[3]);
  assign and_1742_nl = (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1082_nl = (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_697_nl = MUX_s_1_2_2(and_1742_nl, or_1082_nl, MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_1743_nl = (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1081_nl = (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_696_nl = MUX_s_1_2_2(and_1743_nl, or_1081_nl, MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_698_nl = MUX_s_1_2_2(mux_697_nl, mux_696_nl, fsm_output[2]);
  assign and_1744_nl = (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1080_nl = (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_694_nl = MUX_s_1_2_2(and_1744_nl, or_1080_nl, MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_656_nl = ~((~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1078_nl = (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_693_nl = MUX_s_1_2_2(nor_656_nl, or_1078_nl, MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_695_nl = MUX_s_1_2_2(mux_694_nl, mux_693_nl, fsm_output[2]);
  assign mux_699_nl = MUX_s_1_2_2(mux_698_nl, mux_695_nl, fsm_output[3]);
  assign mux_707_nl = MUX_s_1_2_2(mux_706_nl, mux_699_nl, fsm_output[4]);
  assign mux_722_nl = MUX_s_1_2_2(mux_721_nl, mux_707_nl, fsm_output[5]);
  assign and_1745_nl = (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1077_nl = (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_688_nl = MUX_s_1_2_2(and_1745_nl, or_1077_nl, MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_1746_nl = (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1076_nl = (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_687_nl = MUX_s_1_2_2(and_1746_nl, or_1076_nl, MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_689_nl = MUX_s_1_2_2(mux_688_nl, mux_687_nl, fsm_output[2]);
  assign nor_657_nl = ~((~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1074_nl = (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_685_nl = MUX_s_1_2_2(nor_657_nl, or_1074_nl, MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_1747_nl = (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1073_nl = (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_684_nl = MUX_s_1_2_2(and_1747_nl, or_1073_nl, MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_686_nl = MUX_s_1_2_2(mux_685_nl, mux_684_nl, fsm_output[2]);
  assign mux_690_nl = MUX_s_1_2_2(mux_689_nl, mux_686_nl, fsm_output[3]);
  assign nor_658_nl = ~((~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1071_nl = (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_681_nl = MUX_s_1_2_2(nor_658_nl, or_1071_nl, MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_659_nl = ~((~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1069_nl = (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_680_nl = MUX_s_1_2_2(nor_659_nl, or_1069_nl, MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_682_nl = MUX_s_1_2_2(mux_681_nl, mux_680_nl, fsm_output[2]);
  assign nor_660_nl = ~((~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1067_nl = (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_678_nl = MUX_s_1_2_2(nor_660_nl, or_1067_nl, MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_661_nl = ~((~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1065_nl = (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_677_nl = MUX_s_1_2_2(nor_661_nl, or_1065_nl, MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_679_nl = MUX_s_1_2_2(mux_678_nl, mux_677_nl, fsm_output[2]);
  assign mux_683_nl = MUX_s_1_2_2(mux_682_nl, mux_679_nl, fsm_output[3]);
  assign mux_691_nl = MUX_s_1_2_2(mux_690_nl, mux_683_nl, fsm_output[4]);
  assign nor_662_nl = ~((~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1063_nl = (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_673_nl = MUX_s_1_2_2(nor_662_nl, or_1063_nl, MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_663_nl = ~((~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1061_nl = (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_672_nl = MUX_s_1_2_2(nor_663_nl, or_1061_nl, MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_674_nl = MUX_s_1_2_2(mux_673_nl, mux_672_nl, fsm_output[2]);
  assign nor_664_nl = ~((~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1059_nl = (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_670_nl = MUX_s_1_2_2(nor_664_nl, or_1059_nl, MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_665_nl = ~((~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1057_nl = (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_669_nl = MUX_s_1_2_2(nor_665_nl, or_1057_nl, MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_671_nl = MUX_s_1_2_2(mux_670_nl, mux_669_nl, fsm_output[2]);
  assign mux_675_nl = MUX_s_1_2_2(mux_674_nl, mux_671_nl, fsm_output[3]);
  assign nor_666_nl = ~((~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1055_nl = (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_666_nl = MUX_s_1_2_2(nor_666_nl, or_1055_nl, MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nor_667_nl = ~((~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1053_nl = (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_665_nl = MUX_s_1_2_2(nor_667_nl, or_1053_nl, MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_667_nl = MUX_s_1_2_2(mux_666_nl, mux_665_nl, fsm_output[2]);
  assign nor_668_nl = ~((~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]));
  assign or_1051_nl = (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]);
  assign mux_663_nl = MUX_s_1_2_2(nor_668_nl, or_1051_nl, MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign and_1748_nl = (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]);
  assign or_1050_nl = (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7]));
  assign mux_662_nl = MUX_s_1_2_2(and_1748_nl, or_1050_nl, MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_664_nl = MUX_s_1_2_2(mux_663_nl, mux_662_nl, fsm_output[2]);
  assign mux_668_nl = MUX_s_1_2_2(mux_667_nl, mux_664_nl, fsm_output[3]);
  assign mux_676_nl = MUX_s_1_2_2(mux_675_nl, mux_668_nl, fsm_output[4]);
  assign mux_692_nl = MUX_s_1_2_2(mux_691_nl, mux_676_nl, fsm_output[5]);
  assign mux_723_nl = MUX_s_1_2_2(mux_722_nl, mux_692_nl, fsm_output[6]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse = mux_723_nl & and_dcpl_107;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_981;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse = and_dcpl_159 & and_dcpl_1287;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_912;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse = and_dcpl_220 & and_dcpl_1287;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse = and_dcpl_919 & (fsm_output[3])
      & (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & (~ (fsm_output[4])) & nor_225_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse = and_dcpl_159 & and_dcpl_1291;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_922;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse = and_dcpl_220 & and_dcpl_1291;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_928;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse = and_dcpl_159 & and_dcpl_1295;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_933;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse = and_dcpl_220 & and_dcpl_1295;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_939;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse = and_dcpl_159 & and_dcpl_1298;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_944;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse = and_dcpl_220 & and_dcpl_1298;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_949;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse = and_dcpl_159 & and_dcpl_1301;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_953;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse = and_dcpl_220 & and_dcpl_1301;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_958;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse = and_dcpl_159 & and_dcpl_1304;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_962;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse = and_dcpl_220 & and_dcpl_1304;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_966;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse = and_dcpl_159 & and_dcpl_1307;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_970;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse = and_dcpl_220 & and_dcpl_1307;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_974;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse = and_dcpl_1427 & and_dcpl_101;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse = and_dcpl_107 & (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_224 & and_dcpl_162;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse = and_dcpl_1432 & and_dcpl_101;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_981;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse = and_dcpl_1427 & and_dcpl_1287;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_912;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse = and_dcpl_1432 & and_dcpl_1287;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_988;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse = and_dcpl_1427 & and_dcpl_1291;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_922;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse = and_dcpl_1432 & and_dcpl_1291;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_928;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse = and_dcpl_1427 & and_dcpl_1295;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_933;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse = and_dcpl_1432 & and_dcpl_1295;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_939;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse = and_dcpl_1427 & and_dcpl_1298;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse = and_dcpl_1006 & and_dcpl_92
      & (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_943;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse = and_dcpl_1432 & and_dcpl_1298;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_949;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse = and_dcpl_1427 & and_dcpl_1301;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_953;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse = and_dcpl_1432 & and_dcpl_1301;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_958;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse = and_dcpl_1427 & and_dcpl_1304;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_962;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse = and_dcpl_1432 & and_dcpl_1304;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_966;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse = and_dcpl_1427 & and_dcpl_1307;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_970;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse = and_dcpl_1432 & and_dcpl_1307;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_974;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse = and_dcpl_159 & and_dcpl_1326;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1030;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse = and_dcpl_220 & and_dcpl_1326;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1034;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse = and_dcpl_159 & and_dcpl_1329;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1038;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse = and_dcpl_220 & and_dcpl_1329;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1042;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse = and_dcpl_159 & and_dcpl_1332;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1046;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse = and_dcpl_220 & and_dcpl_1332;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1050;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse = and_dcpl_159 & and_dcpl_1335;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1054;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse = and_dcpl_220 & and_dcpl_1335;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1058;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse = and_dcpl_159 & and_dcpl_1338;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1063;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse = and_dcpl_220 & and_dcpl_1338;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse = and_dcpl_919 & (~((MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[4:3]!=2'b00))) & and_1731_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse = and_dcpl_159 & and_dcpl_1341;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse = and_dcpl_108 & and_dcpl_1071
      & (~ (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1731_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse = and_dcpl_220 & and_dcpl_1341;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1075;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse = and_dcpl_159 & and_dcpl_1344;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1079;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse = and_dcpl_220 & and_dcpl_1344;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse = and_dcpl_919 & (~((MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[3]))) & (fsm_output[4]) & and_1731_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse = and_dcpl_159 & and_dcpl_1347;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse = and_dcpl_107 & (~((fsm_output[6])
      | (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))
      & and_dcpl_1087;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse = and_dcpl_220 & and_dcpl_1347;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse = and_dcpl_919 & (fsm_output[3])
      & (~ (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & (fsm_output[4]) & and_1731_cse;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse = and_dcpl_1427 & and_dcpl_1326;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1030;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse = and_dcpl_1432 & and_dcpl_1326;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse = and_dcpl_1101 & (~((MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[4:3]!=2'b00))) & and_dcpl_1029;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse = and_dcpl_1427 & and_dcpl_1329;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1038;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse = and_dcpl_1432 & and_dcpl_1329;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse = and_dcpl_1101 & (fsm_output[3])
      & (~ (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & (~ (fsm_output[4])) & and_dcpl_1029;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse = and_dcpl_1427 & and_dcpl_1332;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1046;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse = and_dcpl_1432 & and_dcpl_1332;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1050;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse = and_dcpl_1427 & and_dcpl_1335;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1054;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse = and_dcpl_1432 & and_dcpl_1335;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1058;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse = and_dcpl_1427 & and_dcpl_1338;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1063;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse = and_dcpl_1432 & and_dcpl_1338;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1125;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse = and_dcpl_1427 & and_dcpl_1341;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1129;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse = and_dcpl_1432 & and_dcpl_1341;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1075;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse = and_dcpl_1427 & and_dcpl_1344;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1079;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse = and_dcpl_1432 & and_dcpl_1344;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1139;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse = and_dcpl_1427 & and_dcpl_1347;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1087;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse = and_dcpl_1432 & and_dcpl_1347;
  assign operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse = and_dcpl_107 & (fsm_output[6])
      & (~ (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_dcpl_1146;
  assign nor_221_cse = ~((fsm_output[1:0]!=2'b00));
  assign or_1557_tmp = ((~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]))
      & (~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_109 & ((~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm)
      | (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva[21]) | (~ MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg)))
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1]))
      & and_dcpl_154);
  assign nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg)}) +
      7'b0000001;
  assign MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1);
  assign MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_ssc = ~(MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_33_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva[21]))
      & MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign nor_250_nl = ~((fsm_output[2]) | and_1698_cse);
  assign mux_213_nl = MUX_s_1_2_2(nor_250_nl, nor_tmp, fsm_output[3]);
  assign and_184_ssc = (~(mux_213_nl | (fsm_output[8]))) & and_dcpl_121;
  assign nor_641_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[5:4]!=2'b00));
  assign nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg)}) +
      7'b0000001;
  assign MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1);
  assign MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_ssc = ~(MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_34_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva[21]))
      & MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_215_nl = MUX_s_1_2_2(not_tmp_273, or_tmp_227, fsm_output[7]);
  assign nor_252_ssc = ~(mux_215_nl | (fsm_output[8]));
  assign nor_616_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[4]));
  assign nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg)}) +
      7'b0000001;
  assign MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1);
  assign MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_ssc = ~(MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_35_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva[21]))
      & MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_217_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_213, fsm_output[7]);
  assign nor_253_ssc = ~(mux_217_nl | (fsm_output[8]));
  assign nor_614_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5);
  assign nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg)}) +
      7'b0000001;
  assign MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1);
  assign MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_ssc = ~(MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_36_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva[21]))
      & MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_219_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_215, fsm_output[7]);
  assign nor_254_ssc = ~(mux_219_nl | (fsm_output[8]));
  assign nor_610_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5);
  assign nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg)}) +
      7'b0000001;
  assign MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1);
  assign MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_ssc = ~(MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_37_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva[21]))
      & MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_221_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_217, fsm_output[7]);
  assign nor_255_ssc = ~(mux_221_nl | (fsm_output[8]));
  assign nor_606_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[4]));
  assign nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg)}) +
      7'b0000001;
  assign MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1);
  assign MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_153_ssc = ~(MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_38_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva[21]))
      & MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_223_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_219, fsm_output[7]);
  assign nor_256_ssc = ~(mux_223_nl | (fsm_output[8]));
  assign nor_600_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[4]));
  assign or_969_cse = (fsm_output[5]) | (fsm_output[7]);
  assign and_1731_cse = (fsm_output[5]) & (fsm_output[7]);
  assign nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg)}) +
      7'b0000001;
  assign MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1);
  assign MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_157_ssc = ~(MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_39_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva[21]))
      & MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_225_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_221, fsm_output[7]);
  assign nor_257_ssc = ~(mux_225_nl | (fsm_output[8]));
  assign nor_598_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5);
  assign nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg)}) +
      7'b0000001;
  assign MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1);
  assign MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_ssc = ~(MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_40_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva[21]))
      & MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_227_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_223, fsm_output[7]);
  assign nor_258_ssc = ~(mux_227_nl | (fsm_output[8]));
  assign nor_594_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[4]));
  assign nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg)}) +
      7'b0000001;
  assign MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1);
  assign MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_165_ssc = ~(MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_41_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva[21]))
      & MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_229_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_225, fsm_output[7]);
  assign nor_259_ssc = ~(mux_229_nl | (fsm_output[8]));
  assign nor_587_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[4]));
  assign or_1164_cse = (fsm_output[2:1]!=2'b00);
  assign nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg)}) +
      7'b0000001;
  assign MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1);
  assign MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_169_ssc = ~(MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_42_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva[21]))
      & MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_231_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_227, fsm_output[7]);
  assign nor_260_ssc = ~(mux_231_nl | (fsm_output[8]));
  assign nor_585_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[4]));
  assign nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg)}) +
      7'b0000001;
  assign MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1);
  assign MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_173_ssc = ~(MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_43_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva[21]))
      & MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_233_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_229, fsm_output[7]);
  assign nor_261_ssc = ~(mux_233_nl | (fsm_output[8]));
  assign nor_581_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5);
  assign nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg)}) +
      7'b0000001;
  assign MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1);
  assign MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_177_ssc = ~(MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_44_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva[21]))
      & MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_234_nl = MUX_s_1_2_2(not_tmp_284, or_dcpl_115, fsm_output[4]);
  assign and_196_ssc = (~ mux_234_nl) & and_dcpl_179;
  assign nor_636_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[5:4]!=2'b00));
  assign nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg)}) +
      7'b0000001;
  assign MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1);
  assign MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_181_ssc = ~(MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_45_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva[21]))
      & MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_236_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_232, fsm_output[7]);
  assign nor_262_ssc = ~(mux_236_nl | (fsm_output[8]));
  assign nor_578_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5);
  assign nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg)}) +
      7'b0000001;
  assign MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1);
  assign MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_185_ssc = ~(MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_46_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva[21]))
      & MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_238_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_234, fsm_output[7]);
  assign nor_263_ssc = ~(mux_238_nl | (fsm_output[8]));
  assign nor_574_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5);
  assign nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg)}) +
      7'b0000001;
  assign MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1);
  assign MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_189_ssc = ~(MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_47_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva[21]))
      & MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_240_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_236, fsm_output[7]);
  assign nor_264_ssc = ~(mux_240_nl | (fsm_output[8]));
  assign nor_568_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[4]));
  assign or_918_cse = (fsm_output[7:6]!=2'b00);
  assign and_1725_cse = (fsm_output[7:6]==2'b11);
  assign nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg)}) +
      7'b0000001;
  assign MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1);
  assign MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_193_ssc = ~(MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_48_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva[21]))
      & MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_242_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_238, fsm_output[7]);
  assign nor_265_ssc = ~(mux_242_nl | (fsm_output[8]));
  assign nor_566_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5);
  assign nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg)}) +
      7'b0000001;
  assign MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1);
  assign MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_197_ssc = ~(MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_49_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva[21]))
      & MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_244_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_240, fsm_output[7]);
  assign nor_266_ssc = ~(mux_244_nl | (fsm_output[8]));
  assign nor_562_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[4]));
  assign nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg)}) +
      7'b0000001;
  assign MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1);
  assign MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_201_ssc = ~(MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_50_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva[21]))
      & MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_246_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_242, fsm_output[7]);
  assign nor_267_ssc = ~(mux_246_nl | (fsm_output[8]));
  assign nor_555_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[4]));
  assign nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg)}) +
      7'b0000001;
  assign MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1);
  assign MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_205_ssc = ~(MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_51_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva[21]))
      & MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_248_nl = MUX_s_1_2_2(not_tmp_273, mux_tmp_244, fsm_output[7]);
  assign nor_268_ssc = ~(mux_248_nl | (fsm_output[8]));
  assign nor_550_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5);
  assign or_1162_cse = nor_550_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6;
  assign nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg)}) +
      7'b0000001;
  assign MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1);
  assign MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_209_ssc = ~(MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_52_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva[21]))
      & MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_249_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_16, fsm_output[7]);
  assign nor_269_ssc = ~(mux_249_nl | (fsm_output[8]));
  assign nor_548_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5);
  assign nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg)}) +
      7'b0000001;
  assign MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1);
  assign MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_213_ssc = ~(MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_53_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva[21]))
      & MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_250_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_17, fsm_output[7]);
  assign nor_270_ssc = ~(mux_250_nl | (fsm_output[8]));
  assign nor_542_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[4]));
  assign or_1161_cse = nor_542_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6;
  assign nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg)}) +
      7'b0000001;
  assign MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1);
  assign MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_217_ssc = ~(MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_54_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva[21]))
      & MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_251_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_18, fsm_output[7]);
  assign nor_271_ssc = ~(mux_251_nl | (fsm_output[8]));
  assign nor_537_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[4]));
  assign or_1160_cse = nor_537_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6;
  assign nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg)}) + 7'b0000001;
  assign MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1);
  assign MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_221_ssc = ~(MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_55_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva[21]))
      & MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_252_nl = MUX_s_1_2_2(not_tmp_284, or_123_cse, fsm_output[4]);
  assign and_210_ssc = (~ mux_252_nl) & and_dcpl_179;
  assign nor_632_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[5:4]!=2'b00));
  assign nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg)}) + 7'b0000001;
  assign MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1);
  assign MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_225_ssc = ~(MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_56_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva[21]))
      & MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_253_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_19, fsm_output[7]);
  assign nor_272_ssc = ~(mux_253_nl | (fsm_output[8]));
  assign nor_533_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[4]));
  assign nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg)}) + 7'b0000001;
  assign MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1);
  assign MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_229_ssc = ~(MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_57_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva[21]))
      & MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_254_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_20, fsm_output[7]);
  assign nor_273_ssc = ~(mux_254_nl | (fsm_output[8]));
  assign nor_528_cse = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[4]));
  assign or_1159_cse = nor_528_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6;
  assign nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg)}) + 7'b0000001;
  assign MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1);
  assign MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_233_ssc = ~(MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_58_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva[21]))
      & MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_255_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_21, fsm_output[7]);
  assign nor_274_ssc = ~(mux_255_nl | (fsm_output[8]));
  assign nor_523_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5);
  assign or_1158_cse = nor_523_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6;
  assign nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg)}) + 7'b0000001;
  assign MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1);
  assign MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_237_ssc = ~(MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_59_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva[21]))
      & MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_256_nl = MUX_s_1_2_2(not_tmp_273, and_tmp_22, fsm_output[7]);
  assign nor_275_ssc = ~(mux_256_nl | (fsm_output[8]));
  assign nor_521_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5);
  assign nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg)}) + 7'b0000001;
  assign MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1);
  assign MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_241_ssc = ~(MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_60_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva[21]))
      & MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_257_nl = MUX_s_1_2_2(not_tmp_284, and_4_cse, fsm_output[4]);
  assign and_219_ssc = (~ mux_257_nl) & and_dcpl_179;
  assign nor_628_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[5:4]!=2'b00));
  assign nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg)}) + 7'b0000001;
  assign MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1);
  assign MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_245_ssc = ~(MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_61_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva[21]))
      & MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign mux_258_nl = MUX_s_1_2_2(not_tmp_284, and_1669_cse, fsm_output[4]);
  assign and_220_ssc = (~ mux_258_nl) & and_dcpl_179;
  assign nor_624_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[5:4]!=2'b00));
  assign nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg)}) + 7'b0000001;
  assign MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1);
  assign MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_249_ssc = ~(MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_62_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva[21]))
      & MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign nor_138_nl = ~((fsm_output[4:2]!=3'b000) | and_1698_cse);
  assign mux_259_nl = MUX_s_1_2_2(nor_138_nl, or_1113_cse, fsm_output[5]);
  assign and_221_ssc = (~ mux_259_nl) & and_dcpl_2;
  assign nor_620_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[5:4]!=2'b00));
  assign nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_s2s_6_7({1'b1 , (~ MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg)}) + 7'b0000001;
  assign MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt
      = nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:0];
  assign nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1);
  assign MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt
      = nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_253_ssc = ~(MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_63_seb
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva[21]))
      & MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign nor_518_cse = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[0])
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4]));
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc = and_dcpl_203 | and_dcpl_154
      | and_dcpl_207;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse = and_dcpl_203 | and_dcpl_154;
  assign ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse = ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse
      & (~ and_dcpl_109);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse
      = and_dcpl_109 | and_dcpl_154;
  assign MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse = ~((z_out_2!=11'b00000000000));
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc = and_dcpl_109
      | and_dcpl_151 | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
      | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_128_nl = ~ MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl
      = MUX_v_11_2_2(11'b00000000000, MAC_ac_float_cctor_m_1_lpi_1_dfm_1, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e1_lt_e2_not_128_nl);
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
      = MUX_v_11_2_2(11'b00000000000, MAC_ac_float_cctor_m_1_lpi_1_dfm_1, MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1);
  assign nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = conv_s2u_11_12(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_nl)
      + conv_s2u_11_12(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl);
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = conv_s2u_11_12(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[11:1])
      + conv_s2u_11_12({result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_10_7
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_6 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_5_4
      , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0});
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm = nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:0];
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0 = $signed((input_m_rsci_idat))
      * $signed((taps_m_rsci_idat[10:0]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0 = $signed(delay_lane_m_33_sva)
      * $signed((taps_m_rsci_idat[373:363]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0 = $signed(delay_lane_m_34_sva)
      * $signed((taps_m_rsci_idat[384:374]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0 = $signed(delay_lane_m_35_sva)
      * $signed((taps_m_rsci_idat[395:385]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0 = $signed(delay_lane_m_36_sva)
      * $signed((taps_m_rsci_idat[406:396]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0 = $signed(delay_lane_m_37_sva)
      * $signed((taps_m_rsci_idat[417:407]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0 = $signed(delay_lane_m_38_sva)
      * $signed((taps_m_rsci_idat[428:418]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0 = $signed(delay_lane_m_39_sva)
      * $signed((taps_m_rsci_idat[439:429]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0 = $signed(delay_lane_m_40_sva)
      * $signed((taps_m_rsci_idat[450:440]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0 = $signed(delay_lane_m_41_sva)
      * $signed((taps_m_rsci_idat[461:451]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0 = $signed(delay_lane_m_42_sva)
      * $signed((taps_m_rsci_idat[472:462]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0 = $signed(delay_lane_m_43_sva)
      * $signed((taps_m_rsci_idat[483:473]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0 = $signed(delay_lane_m_44_sva)
      * $signed((taps_m_rsci_idat[494:484]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0 = $signed(delay_lane_m_45_sva)
      * $signed((taps_m_rsci_idat[505:495]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0 = $signed(delay_lane_m_46_sva)
      * $signed((taps_m_rsci_idat[516:506]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0 = $signed(delay_lane_m_47_sva)
      * $signed((taps_m_rsci_idat[527:517]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0 = $signed(delay_lane_m_48_sva)
      * $signed((taps_m_rsci_idat[538:528]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0 = $signed(delay_lane_m_49_sva)
      * $signed((taps_m_rsci_idat[549:539]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0 = $signed(delay_lane_m_50_sva)
      * $signed((taps_m_rsci_idat[560:550]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0 = $signed(delay_lane_m_51_sva)
      * $signed((taps_m_rsci_idat[571:561]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0 = $signed(delay_lane_m_52_sva)
      * $signed((taps_m_rsci_idat[582:572]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0 = $signed(delay_lane_m_53_sva)
      * $signed((taps_m_rsci_idat[593:583]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0 = $signed(delay_lane_m_54_sva)
      * $signed((taps_m_rsci_idat[604:594]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0 = $signed(delay_lane_m_55_sva)
      * $signed((taps_m_rsci_idat[615:605]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0 = $signed(delay_lane_m_56_sva)
      * $signed((taps_m_rsci_idat[626:616]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0 = $signed(delay_lane_m_57_sva)
      * $signed((taps_m_rsci_idat[637:627]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0 = $signed(delay_lane_m_58_sva)
      * $signed((taps_m_rsci_idat[648:638]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0 = $signed(delay_lane_m_59_sva)
      * $signed((taps_m_rsci_idat[659:649]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0 = $signed(delay_lane_m_60_sva)
      * $signed((taps_m_rsci_idat[670:660]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0 = $signed(delay_lane_m_61_sva)
      * $signed((taps_m_rsci_idat[681:671]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0 = $signed(delay_lane_m_62_sva)
      * $signed((taps_m_rsci_idat[692:682]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0 = $signed(({MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7
      , MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0})) * $signed((taps_m_rsci_idat[703:693]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0 = $signed(delay_lane_m_0_sva)
      * $signed((taps_m_rsci_idat[21:11]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0 = $signed(delay_lane_m_3_sva)
      * $signed((taps_m_rsci_idat[43:33]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0 = $signed(delay_lane_m_4_sva)
      * $signed((taps_m_rsci_idat[54:44]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0 = $signed(delay_lane_m_5_sva)
      * $signed((taps_m_rsci_idat[65:55]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0 = $signed(delay_lane_m_6_sva)
      * $signed((taps_m_rsci_idat[76:66]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0 = $signed(delay_lane_m_7_sva)
      * $signed((taps_m_rsci_idat[87:77]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0 = $signed(delay_lane_m_8_sva)
      * $signed((taps_m_rsci_idat[98:88]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0 = $signed(delay_lane_m_9_sva)
      * $signed((taps_m_rsci_idat[109:99]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0 = $signed(delay_lane_m_10_sva)
      * $signed((taps_m_rsci_idat[120:110]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0 = $signed(delay_lane_m_11_sva)
      * $signed((taps_m_rsci_idat[131:121]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0 = $signed(delay_lane_m_12_sva)
      * $signed((taps_m_rsci_idat[142:132]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0 = $signed(delay_lane_m_13_sva)
      * $signed((taps_m_rsci_idat[153:143]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0 = $signed(delay_lane_m_14_sva)
      * $signed((taps_m_rsci_idat[164:154]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0 = $signed(delay_lane_m_15_sva)
      * $signed((taps_m_rsci_idat[175:165]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0 = $signed(delay_lane_m_16_sva)
      * $signed((taps_m_rsci_idat[186:176]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0 = $signed(delay_lane_m_17_sva)
      * $signed((taps_m_rsci_idat[197:187]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0 = $signed(delay_lane_m_18_sva)
      * $signed((taps_m_rsci_idat[208:198]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0 = $signed(delay_lane_m_19_sva)
      * $signed((taps_m_rsci_idat[219:209]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0 = $signed(delay_lane_m_20_sva)
      * $signed((taps_m_rsci_idat[230:220]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0 = $signed(delay_lane_m_21_sva)
      * $signed((taps_m_rsci_idat[241:231]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0 = $signed(delay_lane_m_22_sva)
      * $signed((taps_m_rsci_idat[252:242]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0 = $signed(delay_lane_m_23_sva)
      * $signed((taps_m_rsci_idat[263:253]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0 = $signed(delay_lane_m_24_sva)
      * $signed((taps_m_rsci_idat[274:264]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0 = $signed(delay_lane_m_25_sva)
      * $signed((taps_m_rsci_idat[285:275]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0 = $signed(delay_lane_m_26_sva)
      * $signed((taps_m_rsci_idat[296:286]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0 = $signed(delay_lane_m_27_sva)
      * $signed((taps_m_rsci_idat[307:297]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0 = $signed(delay_lane_m_28_sva)
      * $signed((taps_m_rsci_idat[318:308]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0 = $signed(delay_lane_m_29_sva)
      * $signed((taps_m_rsci_idat[329:319]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0 = $signed(delay_lane_m_30_sva)
      * $signed((taps_m_rsci_idat[340:330]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0 = $signed(delay_lane_m_31_sva)
      * $signed((taps_m_rsci_idat[351:341]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0 = $signed(delay_lane_m_32_sva)
      * $signed((taps_m_rsci_idat[362:352]));
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0 = $signed(delay_lane_m_1_sva)
      * $signed((taps_m_rsci_idat[32:22]));
  assign nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = conv_s2s_5_6({MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4
      , MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0}) + 6'b000001;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1 = nl_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:0];
  assign MAC_34_r_ac_float_else_and_nl = MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_34_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_34_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_34_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1
      = conv_s2s_6_7({MAC_34_r_ac_float_else_and_nl , MAC_34_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1[6:0];
  assign MAC_35_r_ac_float_else_and_nl = MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_35_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_35_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_35_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1
      = conv_s2s_6_7({MAC_35_r_ac_float_else_and_nl , MAC_35_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1[6:0];
  assign MAC_36_r_ac_float_else_and_nl = MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_36_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_36_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_36_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1
      = conv_s2s_6_7({MAC_36_r_ac_float_else_and_nl , MAC_36_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1[6:0];
  assign MAC_37_r_ac_float_else_and_nl = MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_37_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_37_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_37_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1
      = conv_s2s_6_7({MAC_37_r_ac_float_else_and_nl , MAC_37_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1[6:0];
  assign MAC_38_r_ac_float_else_and_nl = MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_38_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_38_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_38_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1
      = conv_s2s_6_7({MAC_38_r_ac_float_else_and_nl , MAC_38_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1[6:0];
  assign MAC_39_r_ac_float_else_and_nl = MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_39_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_39_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_39_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1
      = conv_s2s_6_7({MAC_39_r_ac_float_else_and_nl , MAC_39_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1[6:0];
  assign MAC_40_r_ac_float_else_and_nl = MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_40_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_40_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_40_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1
      = conv_s2s_6_7({MAC_40_r_ac_float_else_and_nl , MAC_40_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1[6:0];
  assign MAC_41_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5
      & MAC_41_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_41_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0,
      MAC_41_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1
      = conv_s2s_6_7({MAC_41_r_ac_float_else_and_nl , MAC_41_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1[6:0];
  assign MAC_42_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5
      & MAC_42_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_42_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0,
      MAC_42_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1
      = conv_s2s_6_7({MAC_42_r_ac_float_else_and_nl , MAC_42_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1[6:0];
  assign MAC_43_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
      & MAC_43_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_43_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0,
      MAC_43_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1
      = conv_s2s_6_7({MAC_43_r_ac_float_else_and_nl , MAC_43_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1[6:0];
  assign MAC_44_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
      & MAC_44_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_44_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0,
      MAC_44_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1
      = conv_s2s_6_7({MAC_44_r_ac_float_else_and_nl , MAC_44_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1[6:0];
  assign MAC_45_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
      & MAC_45_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_45_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0,
      MAC_45_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1
      = conv_s2s_6_7({MAC_45_r_ac_float_else_and_nl , MAC_45_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1[6:0];
  assign MAC_46_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
      & MAC_46_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_46_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0,
      MAC_46_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1
      = conv_s2s_6_7({MAC_46_r_ac_float_else_and_nl , MAC_46_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1[6:0];
  assign MAC_47_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
      & MAC_47_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_47_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0,
      MAC_47_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1
      = conv_s2s_6_7({MAC_47_r_ac_float_else_and_nl , MAC_47_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1[6:0];
  assign MAC_48_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
      & MAC_48_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_48_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0,
      MAC_48_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1
      = conv_s2s_6_7({MAC_48_r_ac_float_else_and_nl , MAC_48_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1[6:0];
  assign MAC_49_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
      & MAC_49_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_49_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0,
      MAC_49_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1
      = conv_s2s_6_7({MAC_49_r_ac_float_else_and_nl , MAC_49_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1[6:0];
  assign MAC_50_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
      & MAC_50_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_50_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0,
      MAC_50_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1
      = conv_s2s_6_7({MAC_50_r_ac_float_else_and_nl , MAC_50_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1[6:0];
  assign MAC_51_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
      & MAC_51_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_51_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0,
      MAC_51_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1
      = conv_s2s_6_7({MAC_51_r_ac_float_else_and_nl , MAC_51_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1[6:0];
  assign MAC_52_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
      & MAC_52_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_52_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0,
      MAC_52_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1
      = conv_s2s_6_7({MAC_52_r_ac_float_else_and_nl , MAC_52_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1[6:0];
  assign MAC_53_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
      & MAC_53_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_53_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0,
      MAC_53_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1
      = conv_s2s_6_7({MAC_53_r_ac_float_else_and_nl , MAC_53_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1[6:0];
  assign MAC_54_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
      & MAC_54_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_54_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0,
      MAC_54_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1
      = conv_s2s_6_7({MAC_54_r_ac_float_else_and_nl , MAC_54_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1[6:0];
  assign MAC_55_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
      & MAC_55_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_55_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0,
      MAC_55_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1
      = conv_s2s_6_7({MAC_55_r_ac_float_else_and_nl , MAC_55_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1[6:0];
  assign MAC_56_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
      & MAC_56_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_56_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0,
      MAC_56_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1
      = conv_s2s_6_7({MAC_56_r_ac_float_else_and_nl , MAC_56_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1[6:0];
  assign MAC_57_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
      & MAC_57_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_57_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0,
      MAC_57_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1
      = conv_s2s_6_7({MAC_57_r_ac_float_else_and_nl , MAC_57_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1[6:0];
  assign MAC_58_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
      & MAC_58_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_58_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0,
      MAC_58_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1
      = conv_s2s_6_7({MAC_58_r_ac_float_else_and_nl , MAC_58_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1[6:0];
  assign MAC_59_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
      & MAC_59_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_59_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0,
      MAC_59_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1
      = conv_s2s_6_7({MAC_59_r_ac_float_else_and_nl , MAC_59_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1[6:0];
  assign MAC_60_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
      & MAC_60_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_60_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0,
      MAC_60_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1
      = conv_s2s_6_7({MAC_60_r_ac_float_else_and_nl , MAC_60_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1[6:0];
  assign MAC_61_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5
      & MAC_61_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_61_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0,
      MAC_61_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1
      = conv_s2s_6_7({MAC_61_r_ac_float_else_and_nl , MAC_61_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1[6:0];
  assign MAC_62_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
      & MAC_62_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_62_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0,
      MAC_62_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1
      = conv_s2s_6_7({MAC_62_r_ac_float_else_and_nl , MAC_62_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1[6:0];
  assign MAC_63_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
      & MAC_63_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_63_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0,
      MAC_63_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1
      = conv_s2s_6_7({MAC_63_r_ac_float_else_and_nl , MAC_63_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1[6:0];
  assign MAC_1_r_ac_float_else_and_nl = MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_1_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1
      = conv_s2s_6_7({MAC_1_r_ac_float_else_and_nl , MAC_1_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[6:4])
      + 3'b001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign MAC_64_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
      & MAC_64_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_64_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0,
      MAC_64_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1 =
      conv_s2s_6_7({MAC_64_r_ac_float_else_and_nl , MAC_64_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1 = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[10]))
      & MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[10])
      & MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_41_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_162_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_163_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_166_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[10]))
      & MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_167_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[10])
      & MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_42_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_166_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_167_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_170_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[10]))
      & MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_171_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[10])
      & MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_43_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_170_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_171_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_174_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[10]))
      & MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_175_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[10])
      & MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_44_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_174_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_175_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_178_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[10]))
      & MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_179_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[10])
      & MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_45_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_178_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_179_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_182_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[10]))
      & MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_183_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[10])
      & MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_46_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_182_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_183_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_186_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[10]))
      & MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_187_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[10])
      & MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_47_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_186_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_187_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_190_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[10]))
      & MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_191_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[10])
      & MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_48_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_190_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_191_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_194_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[10]))
      & MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_195_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[10])
      & MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_49_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_194_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_195_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0[10]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0[10])
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_18_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_19_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_198_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[10]))
      & MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_199_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[10])
      & MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_50_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_198_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_199_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_202_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[10]))
      & MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_203_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[10])
      & MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_51_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_202_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_203_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_206_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[10]))
      & MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_207_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[10])
      & MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_52_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_206_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_207_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_210_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[10]))
      & MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_211_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[10])
      & MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_53_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_210_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_211_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_214_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[10]))
      & MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_215_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[10])
      & MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_54_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_214_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_215_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_218_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[10]))
      & MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_219_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[10])
      & MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_55_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_218_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_219_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_222_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[10]))
      & MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_223_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[10])
      & MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_56_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_222_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_223_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_226_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[10]))
      & MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_227_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[10])
      & MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_57_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_226_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_227_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_230_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[10]))
      & MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_231_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[10])
      & MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_58_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_230_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_231_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_234_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[10]))
      & MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_235_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[10])
      & MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_59_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_234_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_235_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0[10]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0[10])
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_22_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_23_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_238_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[10]))
      & MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_239_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[10])
      & MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_60_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_238_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_239_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_242_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[10]))
      & MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_243_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[10])
      & MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_61_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_242_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_243_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_246_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[10]))
      & MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_247_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[10])
      & MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_62_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_246_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_247_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_250_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[10]))
      & MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_251_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[10])
      & MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_63_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_250_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_251_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0[10]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0[10])
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_26_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_27_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0[10]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0[10])
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_30_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_31_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0[10])
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_254_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10]))
      & MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_255_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10])
      & MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_254_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_255_nl});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0[10]))
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0[10])
      & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_10_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_11_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      =  -operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1[3:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[1:0]))
      , (~ operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2)}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg)
      + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg)
      + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]))})
      + conv_u2s_5_7(MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)
      + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[4])})
      + 3'b001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg)
      + 7'b0000001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg)
      + 7'b0000001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg)
      + 7'b0000001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg)
      + 7'b0000001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg)
      + 7'b0000001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg)
      + 7'b0000001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg)
      + 7'b0000001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg)
      + 7'b0000001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg)
      + 7'b0000001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg)
      + 7'b0000001;
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[6:4]) + 3'b001;
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp
      = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0[10]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0[10])
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_34_sva_1[3:0];
  assign nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn_oreg) + 7'b0000001;
  assign MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0[10]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0[10])
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_35_sva_1[3:0];
  assign nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn_oreg) + 7'b0000001;
  assign MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0[10]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0[10])
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_36_sva_1[3:0];
  assign nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn_oreg) + 7'b0000001;
  assign MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0[10]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0[10])
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_37_sva_1[3:0];
  assign nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn_oreg) + 7'b0000001;
  assign MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0[10]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0[10])
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_38_sva_1[3:0];
  assign nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn_oreg) + 7'b0000001;
  assign MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0[10]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0[10])
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_39_sva_1[3:0];
  assign nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn_oreg) + 7'b0000001;
  assign MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0[10]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0[10])
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_40_sva_1[3:0];
  assign nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn_oreg) + 7'b0000001;
  assign MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0[10]))
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0[10])
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_41_sva_1[3:0];
  assign nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn_oreg) + 7'b0000001;
  assign MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_lpi_1_dfm_mx0[10]))
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_lpi_1_dfm_mx0[10])
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_42_sva_1[3:0];
  assign nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn_oreg) + 7'b0000001;
  assign MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_lpi_1_dfm_mx0[10]))
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_lpi_1_dfm_mx0[10])
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_43_sva_1[3:0];
  assign nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn_oreg) + 7'b0000001;
  assign MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_lpi_1_dfm_mx0[10]))
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_lpi_1_dfm_mx0[10])
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_44_sva_1[3:0];
  assign nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn_oreg) + 7'b0000001;
  assign MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_lpi_1_dfm_mx0[10]))
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_lpi_1_dfm_mx0[10])
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_45_sva_1[3:0];
  assign nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn_oreg) + 7'b0000001;
  assign MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_lpi_1_dfm_mx0[10]))
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_lpi_1_dfm_mx0[10])
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_46_sva_1[3:0];
  assign nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn_oreg) + 7'b0000001;
  assign MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_lpi_1_dfm_mx0[10]))
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_lpi_1_dfm_mx0[10])
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_47_sva_1[3:0];
  assign nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn_oreg) + 7'b0000001;
  assign MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_lpi_1_dfm_mx0[10]))
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_lpi_1_dfm_mx0[10])
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_48_sva_1[3:0];
  assign nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn_oreg) + 7'b0000001;
  assign MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_lpi_1_dfm_mx0[10]))
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_lpi_1_dfm_mx0[10])
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_25_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_49_sva_1[3:0];
  assign nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn_oreg) + 7'b0000001;
  assign MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_lpi_1_dfm_mx0[10]))
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_lpi_1_dfm_mx0[10])
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_50_sva_1[3:0];
  assign nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn_oreg) + 7'b0000001;
  assign MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_lpi_1_dfm_mx0[10]))
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_lpi_1_dfm_mx0[10])
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_51_sva_1[3:0];
  assign nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn_oreg) + 7'b0000001;
  assign MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_lpi_1_dfm_mx0[10]))
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_lpi_1_dfm_mx0[10])
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_52_sva_1[3:0];
  assign nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn_oreg) + 7'b0000001;
  assign MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_lpi_1_dfm_mx0[10]))
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_lpi_1_dfm_mx0[10])
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_53_sva_1[3:0];
  assign nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn_oreg) + 7'b0000001;
  assign MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_lpi_1_dfm_mx0[10]))
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_lpi_1_dfm_mx0[10])
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_54_sva_1[3:0];
  assign nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn_oreg) + 7'b0000001;
  assign MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_lpi_1_dfm_mx0[10]))
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_lpi_1_dfm_mx0[10])
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_55_sva_1[3:0];
  assign nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn_oreg) + 7'b0000001;
  assign MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_32_lpi_1_dfm_mx0[10]))
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_32_lpi_1_dfm_mx0[10])
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_32_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_32_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_127_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_56_sva_1[3:0];
  assign nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn_oreg) + 7'b0000001;
  assign MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_130_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_33_lpi_1_dfm_mx0[10]))
      & MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_33_lpi_1_dfm_mx0[10])
      & MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_33_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_33_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_130_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_131_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_57_sva_1[3:0];
  assign nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn_oreg) + 7'b0000001;
  assign MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[10]))
      & MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[10])
      & MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_34_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_134_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_135_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_58_sva_1[3:0];
  assign nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn_oreg) + 7'b0000001;
  assign MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_138_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[10]))
      & MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[10])
      & MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_35_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_138_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_139_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_59_sva_1[3:0];
  assign nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn_oreg) + 7'b0000001;
  assign MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_142_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[10]))
      & MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[10])
      & MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_36_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_142_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_143_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_60_sva_1[3:0];
  assign nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn_oreg) + 7'b0000001;
  assign MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_146_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[10]))
      & MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[10])
      & MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_37_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_146_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_147_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_61_sva_1[3:0];
  assign nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn_oreg) + 7'b0000001;
  assign MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_150_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[10]))
      & MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[10])
      & MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_38_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_150_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_151_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_62_sva_1[3:0];
  assign nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn_oreg) + 7'b0000001;
  assign MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_154_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[10]))
      & MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_155_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[10])
      & MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_39_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_154_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_155_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_63_sva_1[3:0];
  assign nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn_oreg) + 7'b0000001;
  assign MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0[10]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0[10])
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w2 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0,
      11'b01111111111, 11'b10000000000, {(~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_14_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_15_nl});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_sva_1[3:0];
  assign nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn_oreg) + 7'b0000001;
  assign MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3 = ~((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[5:4]==2'b01));
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      =  -(MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[3:0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1
      = nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1[3:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_4_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_4_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_5_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_5_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_6_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_6_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_7_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_7_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_8_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_8_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_9_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_9_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_10_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_10_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_11_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_11_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_12_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_12_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_13_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_13_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_14_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_14_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_15_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_15_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_16_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_16_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_17_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_17_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_18_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_18_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_19_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_19_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_20_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_20_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_21_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_21_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_22_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_22_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_23_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_23_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_24_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_24_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_25_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_25_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_26_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_26_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_27_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_27_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_28_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_28_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_29_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_29_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_30_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_30_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_31_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_31_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_32_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_32_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_33_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_33_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1[1]);
  assign MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1])
      | nor_518_cse);
  assign MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6
      | nor_521_cse);
  assign MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6
      | nor_523_cse);
  assign MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6
      | nor_528_cse);
  assign MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
      | nor_533_cse);
  assign MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6
      | nor_537_cse);
  assign MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6
      | nor_542_cse);
  assign MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6
      | nor_548_cse);
  assign MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6
      | nor_550_cse);
  assign MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
      | nor_555_cse);
  assign MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6
      | nor_562_cse);
  assign MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6
      | nor_566_cse);
  assign MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
      | nor_568_cse);
  assign MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6
      | nor_574_cse);
  assign MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6
      | nor_578_cse);
  assign MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6
      | nor_581_cse);
  assign MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6
      | nor_585_cse);
  assign MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
      | nor_587_cse);
  assign MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6
      | nor_594_cse);
  assign MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6
      | nor_598_cse);
  assign MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
      | nor_600_cse);
  assign MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6
      | nor_606_cse);
  assign MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6
      | nor_610_cse);
  assign MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6
      | nor_614_cse);
  assign MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
      | nor_616_cse);
  assign MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6
      | nor_459_cse);
  assign MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6
      | nor_455_cse);
  assign MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6
      | nor_451_cse);
  assign MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
      | nor_447_cse);
  assign MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6
      | nor_442_cse);
  assign MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6
      | nor_438_cse);
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm);
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_32_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_129_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp
      = MUX1HOT_v_7_3_2(MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_32_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_129_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_33_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_64_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm);
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_33_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_33_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm);
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp
      = MUX1HOT_v_7_3_2(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_31_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_125_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_32_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_62_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm);
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_32_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_32_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm);
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp
      = MUX1HOT_v_7_3_2(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_30_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_60_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm);
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm);
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp
      = MUX1HOT_v_7_3_2(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_29_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_58_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm);
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm);
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp
      = MUX1HOT_v_7_3_2(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_28_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_56_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm);
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm);
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp
      = MUX1HOT_v_7_3_2(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_27_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_54_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm);
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm);
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp
      = MUX1HOT_v_7_3_2(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_26_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_52_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm);
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm);
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp
      = MUX1HOT_v_7_3_2(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_25_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_50_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm);
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm);
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp
      = MUX1HOT_v_7_3_2(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_24_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_48_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm);
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp
      = MUX1HOT_v_7_3_2(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_23_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_46_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp
      = MUX1HOT_v_7_3_2(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_22_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_44_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp
      = MUX1HOT_v_7_3_2(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_21_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_42_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp
      = MUX1HOT_v_7_3_2(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_20_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_40_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp
      = MUX1HOT_v_7_3_2(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_19_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_38_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp
      = MUX1HOT_v_7_3_2(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_18_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_36_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp
      = MUX1HOT_v_7_3_2(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_17_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_34_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp
      = MUX1HOT_v_7_3_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_16_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_32_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp
      = MUX1HOT_v_7_3_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_15_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_30_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp
      = MUX1HOT_v_7_3_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_14_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_28_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp
      = MUX1HOT_v_7_3_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_13_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_26_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp
      = MUX1HOT_v_7_3_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_12_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_24_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp
      = MUX1HOT_v_7_3_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_11_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_22_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp
      = MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_10_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_20_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_s2s_6_7({1'b1 , (~ MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp
      = MUX1HOT_v_7_3_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_9_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_18_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp
      = MUX1HOT_v_7_3_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_8_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp
      = MUX1HOT_v_7_3_2(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_7_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_29_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 + conv_u2s_4_7(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp
      = MUX1HOT_v_7_3_2(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_6_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_25_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 + conv_u2s_4_7(result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp
      = MUX1HOT_v_7_3_2(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_5_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_21_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp
      = MUX1HOT_v_7_3_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_4_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_17_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[5:4]!=2'b00))));
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0 + conv_s2s_6_7({1'b1 , (~ MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp
      = MUX1HOT_v_7_3_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_13_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1[1])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm);
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[5:4]!=2'b00))));
  assign or_1042_ssc = MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_cse
      | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0;
  assign MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4 = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1[0])
      & or_1042_ssc;
  assign ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl = ~ or_1042_ssc;
  assign MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0 = MUX_v_4_2_2(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      4'b1111, ac_float_cctor_assign_from_0_0_32_32_AC_TRN_AC_WRAP_if_3_not_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10])
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign MAC_ac_float_cctor_m_1_lpi_1_dfm_1 = MUX1HOT_v_11_3_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva,
      11'b01111111111, 11'b10000000000, {(~ MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1)
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_2_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_3_nl});
  assign nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl = conv_s2s_5_6({(~
      MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_4) , (~ MAC_ac_float_cctor_e_1_lpi_1_dfm_mx0_3_0)})
      + 6'b000001;
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl = nl_MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl[5:0];
  assign MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_itm_5_1 =
      readslicef_6_1_5(MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_nl);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_cse
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1!=2'b00));
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~(operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 | MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4
      = MUX_v_2_2_2(2'b00, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp)
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4!=2'b00))));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_192_mx0
      = MUX_v_4_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm,
      MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_3_lpi_1_dfm_mx0
      = MUX_v_11_2_2((MAC_3_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]),
      (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva + conv_s2s_6_7({1'b1
      , (~ MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0)})
      + 7'b0000001;
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      & (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp
      = MUX1HOT_v_7_3_2(MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      7'b1110000, MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_2_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_9_nl , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_4_tmp,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm);
  assign MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1
      = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[6])
      | (~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[5:4]!=2'b00))));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_195_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_195_nl);
  assign nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = conv_s2s_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      + conv_s2s_5_6({(~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0)
      , (~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1)})
      + 6'b000001;
  assign MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5:0];
  assign MAC_3_result_operator_result_operator_nor_tmp = ~((result_m_1_lpi_1_dfm_1_10_7!=4'b0000)
      | result_m_1_lpi_1_dfm_1_6 | (result_m_1_lpi_1_dfm_1_5_4!=2'b00) | (result_m_1_lpi_1_dfm_1_3_0!=4'b0000));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc
      = ~((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7[3]) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7[3])
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign result_m_1_lpi_1_dfm_1_10_7 = MUX1HOT_v_4_3_2(4'b0111, 4'b1000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7,
      {result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp});
  assign result_m_1_lpi_1_dfm_1_6 = (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc)) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_260_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_318_nl = MUX_v_2_2_2(2'b00,
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_260_nl);
  assign result_m_1_lpi_1_dfm_1_5_4 = MUX_v_2_2_2(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_318_nl,
      2'b11, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_261_nl = ~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_128_ssc;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_319_nl = MUX_v_4_2_2(4'b0000,
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_not_261_nl);
  assign result_m_1_lpi_1_dfm_1_3_0 = MUX_v_4_2_2(result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_319_nl,
      4'b1111, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_64_ssc);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1 = MUX_v_6_2_2(6'b000000,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0);
  assign MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0);
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0);
  assign MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0);
  assign MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0);
  assign MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0);
  assign MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0);
  assign MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0);
  assign MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0);
  assign MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0);
  assign MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0);
  assign MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0);
  assign MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0);
  assign MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0);
  assign MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0);
  assign MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0);
  assign MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0);
  assign MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0);
  assign MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0);
  assign MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0);
  assign MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0);
  assign MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0);
  assign MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0);
  assign MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0);
  assign MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0);
  assign MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0);
  assign MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0);
  assign MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0);
  assign MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0);
  assign MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0);
  assign MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0);
  assign MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp = $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2)
      - $signed(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0);
  assign nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl
      = ({1'b1 , (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva)
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]))})
      + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm)
      + 7'b0000001;
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl
      = nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl[6:0];
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1
      = readslicef_7_1_6(MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_nl);
  assign nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2})
      + conv_s2s_5_6({1'b1 , (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm)})
      + 6'b000001;
  assign MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[5:0];
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp
      = MUX_v_6_2_2(6'b110000, MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_1_itm_6_1);
  assign and_dcpl_1 = ~((fsm_output[8]) | (fsm_output[6]));
  assign and_dcpl_2 = and_dcpl_1 & (~ (fsm_output[7]));
  assign nor_tmp = (fsm_output[2:1]==2'b11);
  assign or_tmp_6 = (fsm_output[4:3]!=2'b00) | nor_tmp;
  assign and_dcpl_10 = ~((fsm_output[8:7]!=2'b00));
  assign or_tmp_49 = (fsm_output[1]) | (fsm_output[6]);
  assign nor_tmp_7 = (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]);
  assign mux_tmp_44 = MUX_s_1_2_2(nor_tmp_7, (fsm_output[6]), fsm_output[3]);
  assign nor_tmp_10 = (fsm_output[3]) & (fsm_output[2]) & (fsm_output[1]) & (fsm_output[6]);
  assign or_tmp_116 = (fsm_output[2]) | (fsm_output[1]) | (fsm_output[6]);
  assign nor_136_cse = ~((fsm_output[3:2]!=2'b00));
  assign or_dcpl_98 = (fsm_output[4:3]!=2'b00) | or_969_cse;
  assign or_dcpl_99 = (fsm_output[6]) | (fsm_output[2]);
  assign or_dcpl_100 = (fsm_output[8]) | (fsm_output[1]);
  assign or_dcpl_103 = or_dcpl_100 | (fsm_output[0]) | or_dcpl_99 | or_dcpl_98;
  assign or_dcpl_105 = (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva)
      | (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[5:4]!=2'b01);
  assign and_dcpl_84 = ~((fsm_output[5:4]!=2'b00));
  assign and_dcpl_85 = and_dcpl_84 & (~ (fsm_output[7]));
  assign and_dcpl_86 = (fsm_output[8]) & (~ (fsm_output[1]));
  assign and_dcpl_92 = ~((fsm_output[4:3]!=2'b00));
  assign and_dcpl_93 = and_dcpl_92 & (~ (fsm_output[5]));
  assign and_dcpl_95 = ~((fsm_output[6]) | (fsm_output[2]));
  assign and_dcpl_97 = and_dcpl_86 & (fsm_output[0]);
  assign and_dcpl_101 = and_dcpl_92 & nor_225_cse;
  assign and_dcpl_102 = ~((fsm_output[8]) | (fsm_output[1]));
  assign and_dcpl_103 = and_dcpl_102 & (~ (fsm_output[0]));
  assign and_dcpl_105 = and_dcpl_103 & and_dcpl_95 & and_dcpl_101;
  assign and_dcpl_106 = (~ (fsm_output[8])) & (fsm_output[1]);
  assign and_dcpl_107 = and_dcpl_106 & (~ (fsm_output[0]));
  assign and_dcpl_108 = and_dcpl_107 & and_dcpl_95;
  assign and_dcpl_109 = and_dcpl_108 & and_dcpl_101;
  assign and_1673_cse = (fsm_output[3:2]==2'b11);
  assign mux_tmp_159 = MUX_s_1_2_2((fsm_output[6]), or_tmp_49, and_1673_cse);
  assign mux_tmp_163 = MUX_s_1_2_2((fsm_output[6]), or_tmp_49, fsm_output[2]);
  assign or_tmp_204 = (fsm_output[5:3]!=3'b000) | mux_tmp_163;
  assign nor_tmp_47 = (fsm_output[4]) & (fsm_output[3]) & (fsm_output[2]) & (fsm_output[6])
      & (fsm_output[1]);
  assign or_tmp_205 = (fsm_output[4]) | (fsm_output[3]) | (fsm_output[2]) | (fsm_output[6])
      | (fsm_output[1]);
  assign nor_tmp_49 = (fsm_output[6]) & (fsm_output[1]);
  assign mux_tmp_166 = MUX_s_1_2_2(nor_tmp_49, (fsm_output[6]), fsm_output[2]);
  assign and_tmp_8 = (fsm_output[4:3]==2'b11) & mux_tmp_166;
  assign and_tmp_9 = (fsm_output[4]) & mux_tmp_44;
  assign and_dcpl_121 = (~((fsm_output[6]) | (fsm_output[4]))) & nor_225_cse;
  assign or_320_nl = (fsm_output[3:2]!=2'b00);
  assign mux_tmp_170 = MUX_s_1_2_2(nor_tmp_49, (fsm_output[6]), or_320_nl);
  assign and_tmp_10 = (fsm_output[4]) & mux_tmp_170;
  assign and_tmp_11 = (fsm_output[3]) & mux_tmp_166;
  assign mux_tmp_172 = MUX_s_1_2_2(and_tmp_11, (fsm_output[6]), fsm_output[4]);
  assign mux_tmp_176 = MUX_s_1_2_2(nor_tmp_49, (fsm_output[6]), or_452_cse);
  assign or_tmp_213 = (fsm_output[1:0]!=2'b10);
  assign or_dcpl_115 = or_1164_cse | (fsm_output[3]);
  assign nor_tmp_53 = (fsm_output[4:1]==4'b1111);
  assign and_tmp_12 = (fsm_output[4:3]==2'b11) & or_1164_cse;
  assign and_tmp_13 = (fsm_output[4]) & or_123_cse;
  assign and_tmp_14 = (fsm_output[4]) & or_dcpl_115;
  assign or_tmp_217 = (fsm_output[4]) | and_1669_cse;
  assign or_tmp_218 = (fsm_output[4]) | and_4_cse;
  assign or_tmp_221 = (fsm_output[3]) | mux_tmp_163;
  assign mux_204_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_221, fsm_output[4]);
  assign or_tmp_222 = (fsm_output[5]) | mux_204_nl;
  assign or_dcpl_120 = (~((fsm_output[8]) & (fsm_output[1]))) | (fsm_output[0]) |
      or_dcpl_99 | or_dcpl_98;
  assign and_dcpl_149 = (~ (fsm_output[6])) & (fsm_output[2]);
  assign and_dcpl_151 = and_dcpl_103 & and_dcpl_149 & and_dcpl_101;
  assign and_dcpl_152 = and_dcpl_106 & (fsm_output[0]);
  assign and_dcpl_153 = and_dcpl_152 & and_dcpl_95;
  assign and_dcpl_154 = and_dcpl_153 & and_dcpl_101;
  assign or_dcpl_126 = or_dcpl_99 | (fsm_output[3]) | or_627_cse | (fsm_output[7]);
  assign and_dcpl_157 = or_dcpl_126 & and_dcpl_152;
  assign and_dcpl_158 = and_dcpl_102 & (fsm_output[0]);
  assign and_dcpl_159 = and_dcpl_158 & and_dcpl_95;
  assign and_dcpl_160 = and_dcpl_159 & and_dcpl_101;
  assign and_dcpl_161 = ~((~((fsm_output[1]) ^ (fsm_output[0]))) | (fsm_output[8]));
  assign and_dcpl_162 = or_dcpl_126 & and_dcpl_161;
  assign or_dcpl_127 = (fsm_output[1:0]!=2'b00);
  assign and_1684_nl = (fsm_output[4:2]==3'b111);
  assign mux_214_nl = MUX_s_1_2_2((fsm_output[6]), or_tmp_49, and_1684_nl);
  assign or_tmp_227 = (fsm_output[5]) | mux_214_nl;
  assign not_tmp_273 = ~((fsm_output[6:2]!=5'b00000) | and_1698_cse);
  assign mux_tmp_213 = MUX_s_1_2_2((fsm_output[6]), or_tmp_205, fsm_output[5]);
  assign or_360_nl = (fsm_output[4:3]!=2'b00) | mux_tmp_163;
  assign mux_tmp_215 = MUX_s_1_2_2((fsm_output[6]), or_360_nl, fsm_output[5]);
  assign or_361_nl = (fsm_output[4]) | mux_80_cse;
  assign mux_tmp_217 = MUX_s_1_2_2((fsm_output[6]), or_361_nl, fsm_output[5]);
  assign or_362_nl = (fsm_output[4]) | mux_tmp_159;
  assign mux_tmp_219 = MUX_s_1_2_2((fsm_output[6]), or_362_nl, fsm_output[5]);
  assign and_1685_cse = (fsm_output[5:4]==2'b11);
  assign mux_tmp_221 = MUX_s_1_2_2((fsm_output[6]), or_224_cse, and_1685_cse);
  assign mux_tmp_223 = MUX_s_1_2_2((fsm_output[6]), or_tmp_221, and_1685_cse);
  assign and_1687_nl = (fsm_output[5:3]==3'b111);
  assign mux_tmp_225 = MUX_s_1_2_2((fsm_output[6]), or_tmp_116, and_1687_nl);
  assign and_1688_nl = (fsm_output[5:2]==4'b1111);
  assign mux_tmp_227 = MUX_s_1_2_2((fsm_output[6]), or_tmp_49, and_1688_nl);
  assign mux_tmp_229 = MUX_s_1_2_2(nor_tmp_49, (fsm_output[6]), or_456_cse);
  assign and_dcpl_179 = and_dcpl_1 & nor_225_cse;
  assign not_tmp_284 = ~((fsm_output[3:2]!=2'b00) | and_1698_cse);
  assign mux_tmp_232 = MUX_s_1_2_2(nor_tmp_7, (fsm_output[6]), or_458_cse);
  assign mux_tmp_234 = MUX_s_1_2_2(and_tmp_11, (fsm_output[6]), or_627_cse);
  assign mux_tmp_236 = MUX_s_1_2_2(nor_tmp_10, (fsm_output[6]), or_627_cse);
  assign mux_tmp_238 = MUX_s_1_2_2(and_tmp_10, (fsm_output[6]), fsm_output[5]);
  assign mux_tmp_240 = MUX_s_1_2_2(and_tmp_9, (fsm_output[6]), fsm_output[5]);
  assign mux_tmp_242 = MUX_s_1_2_2(and_tmp_8, (fsm_output[6]), fsm_output[5]);
  assign mux_tmp_244 = MUX_s_1_2_2(nor_tmp_47, (fsm_output[6]), fsm_output[5]);
  assign and_tmp_16 = (fsm_output[5]) & mux_tmp_176;
  assign and_tmp_17 = (fsm_output[5]) & mux_59_cse;
  assign and_tmp_18 = (fsm_output[5]) & mux_tmp_172;
  assign and_tmp_19 = (fsm_output[5]) & mux_65_cse;
  assign and_tmp_20 = (fsm_output[5:4]==2'b11) & mux_tmp_170;
  assign and_tmp_21 = (fsm_output[5:4]==2'b11) & mux_tmp_44;
  assign and_tmp_22 = (fsm_output[5:3]==3'b111) & mux_tmp_166;
  assign or_dcpl_134 = or_dcpl_100 | (~ (fsm_output[0])) | or_dcpl_99 | or_dcpl_98;
  assign nor_tmp_66 = (fsm_output[6:1]==6'b111111);
  assign and_dcpl_203 = and_dcpl_161 & and_dcpl_95 & and_dcpl_101;
  assign and_dcpl_207 = (fsm_output[8]) & (fsm_output[1]) & (~ (fsm_output[0])) &
      and_dcpl_95 & and_dcpl_101;
  assign and_dcpl_220 = and_dcpl_158 & and_dcpl_149;
  assign and_dcpl_221 = and_dcpl_220 & and_dcpl_101;
  assign and_dcpl_223 = nor_136_cse & (~ (fsm_output[4]));
  assign and_dcpl_224 = and_dcpl_223 & nor_225_cse;
  assign and_dcpl_225 = ~((fsm_output[6]) | (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_dcpl_235 = ~((fsm_output[6]) | (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign mux_264_nl = MUX_s_1_2_2((~ (fsm_output[8])), (fsm_output[8]), fsm_output[6]);
  assign or_391_nl = (~ (fsm_output[6])) | (fsm_output[8]);
  assign mux_265_nl = MUX_s_1_2_2(mux_264_nl, or_391_nl, fsm_output[2]);
  assign mux_266_nl = MUX_s_1_2_2(mux_265_nl, (fsm_output[8]), or_150_cse);
  assign and_dcpl_245 = (~ mux_266_nl) & nor_221_cse;
  assign and_dcpl_259 = and_dcpl_95 & (~ (fsm_output[3]));
  assign and_dcpl_260 = and_dcpl_107 & and_dcpl_259;
  assign or_dcpl_150 = or_152_cse | (fsm_output[7]);
  assign and_dcpl_497 = and_dcpl_259 & and_dcpl_85;
  assign or_dcpl_172 = (fsm_output[8:7]!=2'b00);
  assign mux_tmp_294 = MUX_s_1_2_2((~ (fsm_output[1])), (fsm_output[1]), fsm_output[6]);
  assign or_tmp_285 = (fsm_output[6]) | (~ or_tmp_213);
  assign and_dcpl_546 = and_dcpl_149 & (~ (fsm_output[3]));
  assign and_dcpl_547 = and_dcpl_546 & and_dcpl_85;
  assign mux_tmp_314 = MUX_s_1_2_2((~ (fsm_output[1])), (fsm_output[1]), fsm_output[0]);
  assign or_tmp_292 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign or_tmp_297 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_308 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_314 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_318 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_326 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_330 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_334 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_346 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_356 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_362 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_370 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_tmp_374 = (fsm_output[7]) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign and_dcpl_556 = and_dcpl_95 & (fsm_output[3]);
  assign and_dcpl_561 = and_dcpl_149 & (fsm_output[3]);
  assign and_dcpl_566 = (fsm_output[5:4]==2'b01);
  assign and_dcpl_567 = and_dcpl_566 & (~ (fsm_output[7]));
  assign and_dcpl_584 = (fsm_output[5:4]==2'b10);
  assign and_dcpl_585 = and_dcpl_584 & (~ (fsm_output[7]));
  assign and_dcpl_603 = and_1685_cse & (~ (fsm_output[7]));
  assign and_dcpl_620 = (fsm_output[6]) & (~ (fsm_output[2]));
  assign and_dcpl_621 = and_dcpl_620 & (~ (fsm_output[3]));
  assign and_dcpl_626 = (fsm_output[6]) & (fsm_output[2]);
  assign and_dcpl_627 = and_dcpl_626 & (~ (fsm_output[3]));
  assign and_dcpl_632 = and_dcpl_620 & (fsm_output[3]);
  assign and_dcpl_637 = and_dcpl_626 & (fsm_output[3]);
  assign and_dcpl_690 = and_dcpl_84 & (fsm_output[7]);
  assign and_dcpl_707 = and_dcpl_566 & (fsm_output[7]);
  assign and_dcpl_724 = and_dcpl_584 & (fsm_output[7]);
  assign and_dcpl_741 = and_1685_cse & (fsm_output[7]);
  assign or_dcpl_278 = or_152_cse | (fsm_output[4]) | or_969_cse;
  assign not_tmp_640 = ~((fsm_output[6:2]!=5'b00000));
  assign or_1133_cse = (fsm_output[6:4]!=3'b000);
  assign nor_tmp_76 = or_1133_cse & (fsm_output[7]);
  assign mux_tmp_468 = MUX_s_1_2_2((~ (fsm_output[7])), (fsm_output[7]), or_1133_cse);
  assign or_dcpl_308 = (fsm_output[6]) | (fsm_output[3]) | (fsm_output[4]) | or_969_cse;
  assign and_dcpl_910 = (fsm_output[3:2]==2'b10);
  assign and_dcpl_911 = and_dcpl_910 & (~ (fsm_output[4]));
  assign and_dcpl_912 = and_dcpl_911 & nor_225_cse;
  assign and_dcpl_919 = and_dcpl_107 & and_dcpl_149;
  assign and_dcpl_921 = nor_136_cse & (fsm_output[4]);
  assign and_dcpl_922 = and_dcpl_921 & nor_225_cse;
  assign and_dcpl_926 = (fsm_output[3:2]==2'b01);
  assign and_dcpl_927 = and_dcpl_926 & (fsm_output[4]);
  assign and_dcpl_928 = and_dcpl_927 & nor_225_cse;
  assign and_dcpl_932 = and_dcpl_910 & (fsm_output[4]);
  assign and_dcpl_933 = and_dcpl_932 & nor_225_cse;
  assign and_dcpl_938 = and_1673_cse & (fsm_output[4]);
  assign and_dcpl_939 = and_dcpl_938 & nor_225_cse;
  assign and_dcpl_943 = (fsm_output[5]) & (~ (fsm_output[7]));
  assign and_dcpl_944 = and_dcpl_223 & and_dcpl_943;
  assign and_dcpl_948 = and_dcpl_926 & (~ (fsm_output[4]));
  assign and_dcpl_949 = and_dcpl_948 & and_dcpl_943;
  assign and_dcpl_953 = and_dcpl_911 & and_dcpl_943;
  assign and_dcpl_957 = and_1673_cse & (~ (fsm_output[4]));
  assign and_dcpl_958 = and_dcpl_957 & and_dcpl_943;
  assign and_dcpl_962 = and_dcpl_921 & and_dcpl_943;
  assign and_dcpl_966 = and_dcpl_927 & and_dcpl_943;
  assign and_dcpl_970 = and_dcpl_932 & and_dcpl_943;
  assign and_dcpl_974 = and_dcpl_938 & and_dcpl_943;
  assign and_dcpl_981 = and_dcpl_948 & nor_225_cse;
  assign and_dcpl_988 = and_dcpl_957 & nor_225_cse;
  assign and_dcpl_1006 = and_dcpl_107 & and_dcpl_620;
  assign and_dcpl_1029 = (~ (fsm_output[5])) & (fsm_output[7]);
  assign and_dcpl_1030 = and_dcpl_223 & and_dcpl_1029;
  assign and_dcpl_1034 = and_dcpl_948 & and_dcpl_1029;
  assign and_dcpl_1038 = and_dcpl_911 & and_dcpl_1029;
  assign and_dcpl_1042 = and_dcpl_957 & and_dcpl_1029;
  assign and_dcpl_1046 = and_dcpl_921 & and_dcpl_1029;
  assign and_dcpl_1050 = and_dcpl_927 & and_dcpl_1029;
  assign and_dcpl_1054 = and_dcpl_932 & and_dcpl_1029;
  assign and_dcpl_1058 = and_dcpl_938 & and_dcpl_1029;
  assign and_dcpl_1063 = and_dcpl_223 & and_1731_cse;
  assign and_dcpl_1071 = (fsm_output[4:3]==2'b01);
  assign and_dcpl_1075 = and_dcpl_957 & and_1731_cse;
  assign and_dcpl_1079 = and_dcpl_921 & and_1731_cse;
  assign and_dcpl_1087 = and_dcpl_932 & and_1731_cse;
  assign and_dcpl_1101 = and_dcpl_107 & and_dcpl_626;
  assign and_dcpl_1125 = and_dcpl_948 & and_1731_cse;
  assign and_dcpl_1129 = and_dcpl_911 & and_1731_cse;
  assign and_dcpl_1139 = and_dcpl_927 & and_1731_cse;
  assign and_dcpl_1146 = and_dcpl_938 & and_1731_cse;
  assign and_1695_cse = (fsm_output[7:3]==5'b11111);
  assign or_dcpl_316 = (~ (fsm_output[1])) | (fsm_output[8]) | (~ (fsm_output[0]))
      | or_dcpl_99 | or_dcpl_98;
  assign nor_246_nl = ~((fsm_output[7:4]!=4'b0000));
  assign and_1697_nl = (fsm_output[7:4]==4'b1111);
  assign mux_tmp_557 = MUX_s_1_2_2(nor_246_nl, and_1697_nl, fsm_output[3]);
  assign or_tmp_589 = (fsm_output[5:1]!=5'b00000);
  assign or_dcpl_368 = or_152_cse | or_969_cse;
  assign and_dcpl_1276 = (fsm_output[1:0]==2'b01);
  assign and_dcpl_1287 = and_dcpl_1071 & nor_225_cse;
  assign and_dcpl_1290 = (fsm_output[4:3]==2'b10);
  assign and_dcpl_1291 = and_dcpl_1290 & nor_225_cse;
  assign and_dcpl_1295 = and_1670_cse & nor_225_cse;
  assign and_dcpl_1298 = and_dcpl_92 & and_dcpl_943;
  assign and_dcpl_1301 = and_dcpl_1071 & and_dcpl_943;
  assign and_dcpl_1304 = and_dcpl_1290 & and_dcpl_943;
  assign and_dcpl_1307 = and_1670_cse & and_dcpl_943;
  assign and_dcpl_1326 = and_dcpl_92 & and_dcpl_1029;
  assign and_dcpl_1329 = and_dcpl_1071 & and_dcpl_1029;
  assign and_dcpl_1332 = and_dcpl_1290 & and_dcpl_1029;
  assign and_dcpl_1335 = and_1670_cse & and_dcpl_1029;
  assign and_dcpl_1338 = and_dcpl_92 & and_1731_cse;
  assign and_dcpl_1341 = and_dcpl_1071 & and_1731_cse;
  assign and_dcpl_1344 = and_dcpl_1290 & and_1731_cse;
  assign and_dcpl_1347 = and_1670_cse & and_1731_cse;
  assign and_dcpl_1427 = and_dcpl_158 & and_dcpl_620;
  assign and_dcpl_1432 = and_dcpl_158 & and_dcpl_626;
  assign return_e_rsci_idat_mx0c1 = and_dcpl_97 & and_dcpl_95 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      & and_dcpl_93 & (~((fsm_output[7]) | (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[5])))
      & (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[4]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 = or_dcpl_127
      & (~ (fsm_output[8])) & and_dcpl_95 & and_dcpl_101;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
      = and_dcpl_153 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
      = and_dcpl_153 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c0
      = and_dcpl_107 & (~ (fsm_output[6])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2])
      & and_dcpl_224;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c1
      = and_dcpl_107 & (~((fsm_output[6]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2])))
      & and_dcpl_224;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c0
      = and_dcpl_107 & (~ (fsm_output[6])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2])
      & and_dcpl_224;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c1
      = and_dcpl_107 & (~((fsm_output[6]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2])))
      & and_dcpl_224;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
      = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
      = and_dcpl_108 & and_dcpl_93 & (~((fsm_output[7]) | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3 = or_dcpl_308
      & and_dcpl_158;
  assign or_1135_nl = (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_486_nl = ~((MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_546_nl = MUX_s_1_2_2(or_1135_nl, nor_486_nl, MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_547_nl = MUX_s_1_2_2(nor_369_cse, mux_546_nl, fsm_output[2]);
  assign or_1136_nl = (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_487_nl = ~((MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_544_nl = MUX_s_1_2_2(or_1136_nl, nor_487_nl, MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1137_nl = (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_488_nl = ~((MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_543_nl = MUX_s_1_2_2(or_1137_nl, nor_488_nl, MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_545_nl = MUX_s_1_2_2(mux_544_nl, mux_543_nl, fsm_output[2]);
  assign mux_548_nl = MUX_s_1_2_2(mux_547_nl, mux_545_nl, fsm_output[3]);
  assign or_1138_nl = (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_489_nl = ~((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_540_nl = MUX_s_1_2_2(or_1138_nl, nor_489_nl, MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1139_nl = (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_490_nl = ~((MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_539_nl = MUX_s_1_2_2(or_1139_nl, nor_490_nl, MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_541_nl = MUX_s_1_2_2(mux_540_nl, mux_539_nl, fsm_output[2]);
  assign or_1140_nl = (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_491_nl = ~((MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_537_nl = MUX_s_1_2_2(or_1140_nl, nor_491_nl, MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1141_nl = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_492_nl = ~((MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_536_nl = MUX_s_1_2_2(or_1141_nl, nor_492_nl, MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_538_nl = MUX_s_1_2_2(mux_537_nl, mux_536_nl, fsm_output[2]);
  assign mux_542_nl = MUX_s_1_2_2(mux_541_nl, mux_538_nl, fsm_output[3]);
  assign mux_549_nl = MUX_s_1_2_2(mux_548_nl, mux_542_nl, fsm_output[4]);
  assign or_1142_nl = (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_493_nl = ~((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_532_nl = MUX_s_1_2_2(or_1142_nl, nor_493_nl, MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nand_47_nl = ~((MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_494_nl = ~((MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_531_nl = MUX_s_1_2_2(nand_47_nl, nor_494_nl, MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_533_nl = MUX_s_1_2_2(mux_532_nl, mux_531_nl, fsm_output[2]);
  assign or_1143_nl = (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_495_nl = ~((MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_529_nl = MUX_s_1_2_2(or_1143_nl, nor_495_nl, MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1144_nl = (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_496_nl = ~((MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_528_nl = MUX_s_1_2_2(or_1144_nl, nor_496_nl, MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_530_nl = MUX_s_1_2_2(mux_529_nl, mux_528_nl, fsm_output[2]);
  assign mux_534_nl = MUX_s_1_2_2(mux_533_nl, mux_530_nl, fsm_output[3]);
  assign nand_48_nl = ~((MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_497_nl = ~((MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_525_nl = MUX_s_1_2_2(nand_48_nl, nor_497_nl, MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nand_49_nl = ~((MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_498_nl = ~((MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_524_nl = MUX_s_1_2_2(nand_49_nl, nor_498_nl, MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_526_nl = MUX_s_1_2_2(mux_525_nl, mux_524_nl, fsm_output[2]);
  assign nand_50_nl = ~((MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_499_nl = ~((MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_522_nl = MUX_s_1_2_2(nand_50_nl, nor_499_nl, MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1145_nl = (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_500_nl = ~((MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_521_nl = MUX_s_1_2_2(or_1145_nl, nor_500_nl, MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_523_nl = MUX_s_1_2_2(mux_522_nl, mux_521_nl, fsm_output[2]);
  assign mux_527_nl = MUX_s_1_2_2(mux_526_nl, mux_523_nl, fsm_output[3]);
  assign mux_535_nl = MUX_s_1_2_2(mux_534_nl, mux_527_nl, fsm_output[4]);
  assign mux_550_nl = MUX_s_1_2_2(mux_549_nl, mux_535_nl, fsm_output[5]);
  assign nand_51_nl = ~((MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_501_nl = ~((MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_516_nl = MUX_s_1_2_2(nand_51_nl, nor_501_nl, MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nand_52_nl = ~((MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_502_nl = ~((MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_515_nl = MUX_s_1_2_2(nand_52_nl, nor_502_nl, MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_517_nl = MUX_s_1_2_2(mux_516_nl, mux_515_nl, fsm_output[2]);
  assign or_1146_nl = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_503_nl = ~((MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_513_nl = MUX_s_1_2_2(or_1146_nl, nor_503_nl, MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nand_53_nl = ~((MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_504_nl = ~((MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_512_nl = MUX_s_1_2_2(nand_53_nl, nor_504_nl, MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_514_nl = MUX_s_1_2_2(mux_513_nl, mux_512_nl, fsm_output[2]);
  assign mux_518_nl = MUX_s_1_2_2(mux_517_nl, mux_514_nl, fsm_output[3]);
  assign or_1147_nl = (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_505_nl = ~((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_509_nl = MUX_s_1_2_2(or_1147_nl, nor_505_nl, MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1148_nl = (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_506_nl = ~((MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_508_nl = MUX_s_1_2_2(or_1148_nl, nor_506_nl, MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_510_nl = MUX_s_1_2_2(mux_509_nl, mux_508_nl, fsm_output[2]);
  assign or_1149_nl = (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_507_nl = ~((MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_506_nl = MUX_s_1_2_2(or_1149_nl, nor_507_nl, MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1150_nl = (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_508_nl = ~((MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_505_nl = MUX_s_1_2_2(or_1150_nl, nor_508_nl, MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_507_nl = MUX_s_1_2_2(mux_506_nl, mux_505_nl, fsm_output[2]);
  assign mux_511_nl = MUX_s_1_2_2(mux_510_nl, mux_507_nl, fsm_output[3]);
  assign mux_519_nl = MUX_s_1_2_2(mux_518_nl, mux_511_nl, fsm_output[4]);
  assign or_1151_nl = (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_509_nl = ~((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_501_nl = MUX_s_1_2_2(or_1151_nl, nor_509_nl, MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1152_nl = (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_510_nl = ~((MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_500_nl = MUX_s_1_2_2(or_1152_nl, nor_510_nl, MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_502_nl = MUX_s_1_2_2(mux_501_nl, mux_500_nl, fsm_output[2]);
  assign or_1153_nl = (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_511_nl = ~((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_498_nl = MUX_s_1_2_2(or_1153_nl, nor_511_nl, MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1154_nl = (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_512_nl = ~((MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_497_nl = MUX_s_1_2_2(or_1154_nl, nor_512_nl, MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_499_nl = MUX_s_1_2_2(mux_498_nl, mux_497_nl, fsm_output[2]);
  assign mux_503_nl = MUX_s_1_2_2(mux_502_nl, mux_499_nl, fsm_output[3]);
  assign or_1155_nl = (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_513_nl = ~((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_494_nl = MUX_s_1_2_2(or_1155_nl, nor_513_nl, MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign or_1156_nl = (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_514_nl = ~((MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_493_nl = MUX_s_1_2_2(or_1156_nl, nor_514_nl, MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_495_nl = MUX_s_1_2_2(mux_494_nl, mux_493_nl, fsm_output[2]);
  assign or_1157_nl = (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      | (fsm_output[7]);
  assign nor_515_nl = ~((MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (fsm_output[7]));
  assign mux_491_nl = MUX_s_1_2_2(or_1157_nl, nor_515_nl, MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign nand_54_nl = ~((MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[7]));
  assign nor_516_nl = ~((MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      | (~ (fsm_output[7])));
  assign mux_490_nl = MUX_s_1_2_2(nand_54_nl, nor_516_nl, MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_492_nl = MUX_s_1_2_2(mux_491_nl, mux_490_nl, fsm_output[2]);
  assign mux_496_nl = MUX_s_1_2_2(mux_495_nl, mux_492_nl, fsm_output[3]);
  assign mux_504_nl = MUX_s_1_2_2(mux_503_nl, mux_496_nl, fsm_output[4]);
  assign mux_520_nl = MUX_s_1_2_2(mux_519_nl, mux_504_nl, fsm_output[5]);
  assign mux_551_nl = MUX_s_1_2_2(mux_550_nl, mux_520_nl, fsm_output[6]);
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
      = mux_551_nl & and_dcpl_107;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_912;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
      = and_dcpl_919 & (fsm_output[3]) & (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ (fsm_output[4])) & nor_225_cse;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_922;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_928;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_933;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_939;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_944;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_949;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_953;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_958;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_962;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_966;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_970;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_974;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
      = and_dcpl_107 & (fsm_output[6]) & (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_224;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
      = and_dcpl_107 & (fsm_output[6]) & (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_981;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
      = and_dcpl_107 & (fsm_output[6]) & (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_912;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
      = and_dcpl_107 & (fsm_output[6]) & (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_988;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
      = and_dcpl_107 & (fsm_output[6]) & (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_922;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
      = and_dcpl_107 & (fsm_output[6]) & (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_928;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
      = and_dcpl_107 & (fsm_output[6]) & (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_933;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
      = and_dcpl_107 & (fsm_output[6]) & (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_939;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
      = and_dcpl_1006 & and_dcpl_92 & (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_943;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
      = and_dcpl_107 & (fsm_output[6]) & (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_949;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
      = and_dcpl_107 & (fsm_output[6]) & (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_953;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
      = and_dcpl_107 & (fsm_output[6]) & (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_958;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
      = and_dcpl_107 & (fsm_output[6]) & (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_962;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
      = and_dcpl_107 & (fsm_output[6]) & (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_966;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
      = and_dcpl_107 & (fsm_output[6]) & (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_970;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
      = and_dcpl_107 & (fsm_output[6]) & (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_974;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1030;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1034;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1038;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1042;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1046;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1050;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1054;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1058;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1063;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
      = and_dcpl_919 & (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[4:3]==2'b00) & and_1731_cse;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
      = and_dcpl_108 & and_dcpl_1071 & (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1731_cse;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1075;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1079;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
      = and_dcpl_919 & (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[4:3]==2'b10) & and_1731_cse;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
      = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1087;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
      = and_dcpl_919 & (fsm_output[3]) & (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[4]) & and_1731_cse;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
      = and_dcpl_107 & (fsm_output[6]) & (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1030;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
      = and_dcpl_1101 & (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (fsm_output[4:3]==2'b00) & and_dcpl_1029;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
      = and_dcpl_107 & (fsm_output[6]) & (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1038;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
      = and_dcpl_1101 & (fsm_output[3]) & (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ (fsm_output[4])) & and_dcpl_1029;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
      = and_dcpl_107 & (fsm_output[6]) & (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1046;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
      = and_dcpl_107 & (fsm_output[6]) & (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1050;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
      = and_dcpl_107 & (fsm_output[6]) & (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1054;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
      = and_dcpl_107 & (fsm_output[6]) & (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1058;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
      = and_dcpl_107 & (fsm_output[6]) & (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1063;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
      = and_dcpl_107 & (fsm_output[6]) & (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1125;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
      = and_dcpl_107 & (fsm_output[6]) & (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1129;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
      = and_dcpl_107 & (fsm_output[6]) & (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1075;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
      = and_dcpl_107 & (fsm_output[6]) & (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1079;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
      = and_dcpl_107 & (fsm_output[6]) & (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1139;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
      = and_dcpl_107 & (fsm_output[6]) & (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1087;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64
      = and_dcpl_107 & (fsm_output[6]) & (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_dcpl_1146;
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]))})
      + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg) + 7'b0000001;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg)
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg)
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg)
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg)
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg)
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg)
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg)
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg)
      + 7'b0000001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg)
      + 7'b0000001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg)
      + 7'b0000001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg)
      + 7'b0000001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg)
      + 7'b0000001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg)
      + 7'b0000001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg)
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg)
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg)
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg)
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg)
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = ({1'b1 , (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[1:0]))
      , (~ (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]))}) + conv_u2s_5_7(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg)
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl[6:0];
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      = readslicef_7_1_6(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_nl);
  assign or_tmp_717 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm;
  assign or_tmp_718 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm;
  assign or_tmp_719 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm;
  assign or_tmp_725 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  assign or_tmp_731 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva;
  assign or_tmp_734 = and_dcpl_1301 | and_dcpl_1347;
  assign mux_tmp = MUX_s_1_2_2(and_dcpl_1301, or_tmp_734, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign nor_tmp_132 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
      & and_dcpl_1347;
  assign mux_724_nl = MUX_s_1_2_2(nor_tmp_132, mux_tmp, or_tmp_731);
  assign or_1188_nl = (or_tmp_731 & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_722 = MUX_s_1_2_2(mux_724_nl, or_1188_nl, ac_float_cctor_operator_return_sva);
  assign or_1191_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | mux_tmp_722;
  assign mux_tmp_723 = MUX_s_1_2_2(mux_tmp_722, or_1191_nl, and_dcpl_1295);
  assign or_1192_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_723;
  assign mux_tmp_724 = MUX_s_1_2_2(mux_tmp_723, or_1192_nl, and_dcpl_1332);
  assign or_1193_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | mux_tmp_724;
  assign mux_tmp_725 = MUX_s_1_2_2(mux_tmp_724, or_1193_nl, and_dcpl_1304);
  assign or_1194_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | mux_tmp_725;
  assign mux_tmp_726 = MUX_s_1_2_2(mux_tmp_725, or_1194_nl, and_dcpl_1291);
  assign or_1195_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | mux_tmp_726;
  assign mux_tmp_727 = MUX_s_1_2_2(mux_tmp_726, or_1195_nl, and_dcpl_1307);
  assign or_1196_nl = or_tmp_725 | mux_tmp_727;
  assign mux_tmp_728 = MUX_s_1_2_2(mux_tmp_727, or_1196_nl, and_dcpl_101);
  assign or_1197_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_728;
  assign mux_tmp_729 = MUX_s_1_2_2(mux_tmp_728, or_1197_nl, and_dcpl_1287);
  assign or_1198_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | mux_tmp_729;
  assign mux_tmp_730 = MUX_s_1_2_2(mux_tmp_729, or_1198_nl, and_dcpl_1298);
  assign or_1199_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_730;
  assign mux_tmp_731 = MUX_s_1_2_2(mux_tmp_730, or_1199_nl, and_dcpl_1338);
  assign or_1200_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | mux_tmp_731;
  assign mux_tmp_732 = MUX_s_1_2_2(mux_tmp_731, or_1200_nl, and_dcpl_1344);
  assign or_tmp_746 = and_dcpl_919 | and_dcpl_108;
  assign or_tmp_747 = or_tmp_746 | mux_tmp_732;
  assign or_1201_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
      | and_dcpl_919 | and_dcpl_108 | mux_tmp_732;
  assign mux_tmp_733 = MUX_s_1_2_2(or_tmp_747, or_1201_nl, and_dcpl_1335);
  assign or_tmp_748 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm;
  assign or_tmp_762 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm;
  assign mux_tmp_734 = MUX_s_1_2_2(and_dcpl_1301, or_tmp_734, or_tmp_762);
  assign mux_tmp_735 = MUX_s_1_2_2(and_dcpl_1301, or_tmp_734, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm);
  assign nor_tmp_135 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm
      & and_dcpl_1347;
  assign mux_tmp_736 = MUX_s_1_2_2(nor_tmp_135, mux_tmp_735, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva);
  assign or_1219_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_737 = MUX_s_1_2_2(mux_tmp_736, or_1219_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign mux_741_nl = MUX_s_1_2_2(mux_tmp_737, mux_tmp_734, or_tmp_731);
  assign or_1216_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva)
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_739 = MUX_s_1_2_2(mux_741_nl, or_1216_nl, ac_float_cctor_operator_return_sva);
  assign or_1220_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_739;
  assign mux_tmp_740 = MUX_s_1_2_2(mux_tmp_739, or_1220_nl, and_dcpl_1295);
  assign or_1221_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_740;
  assign mux_tmp_741 = MUX_s_1_2_2(mux_tmp_740, or_1221_nl, and_dcpl_1332);
  assign or_1222_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_741;
  assign mux_tmp_742 = MUX_s_1_2_2(mux_tmp_741, or_1222_nl, and_dcpl_1304);
  assign or_1223_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | mux_tmp_742;
  assign mux_tmp_743 = MUX_s_1_2_2(mux_tmp_742, or_1223_nl, and_dcpl_1291);
  assign or_1224_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_743;
  assign mux_tmp_744 = MUX_s_1_2_2(mux_tmp_743, or_1224_nl, and_dcpl_1307);
  assign or_1225_nl = or_tmp_725 | mux_tmp_744;
  assign mux_tmp_745 = MUX_s_1_2_2(mux_tmp_744, or_1225_nl, and_dcpl_101);
  assign or_1226_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_745;
  assign mux_tmp_746 = MUX_s_1_2_2(mux_tmp_745, or_1226_nl, and_dcpl_1287);
  assign or_1227_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_746;
  assign mux_tmp_747 = MUX_s_1_2_2(mux_tmp_746, or_1227_nl, and_dcpl_1298);
  assign or_1228_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_747;
  assign mux_tmp_748 = MUX_s_1_2_2(mux_tmp_747, or_1228_nl, and_dcpl_1338);
  assign or_1229_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | mux_tmp_748;
  assign mux_752_nl = MUX_s_1_2_2(mux_tmp_748, or_1229_nl, and_dcpl_1344);
  assign mux_tmp_750 = MUX_s_1_2_2(mux_tmp_732, mux_752_nl, and_dcpl_108);
  assign or_tmp_774 = and_dcpl_919 | mux_tmp_750;
  assign mux_tmp_751 = MUX_s_1_2_2(or_tmp_774, or_tmp_747, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign or_1231_nl = or_tmp_748 | mux_tmp_751;
  assign mux_tmp_752 = MUX_s_1_2_2(or_tmp_774, or_1231_nl, and_dcpl_1335);
  assign or_tmp_776 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva;
  assign or_tmp_777 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm;
  assign or_tmp_783 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  assign nor_tmp_137 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm
      & and_dcpl_1347;
  assign or_tmp_792 = and_dcpl_1301 | nor_tmp_137;
  assign mux_tmp_754 = MUX_s_1_2_2(or_tmp_792, or_tmp_734, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign and_1766_cse = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      & and_dcpl_1301;
  assign or_tmp_793 = and_1766_cse | and_dcpl_1347;
  assign or_tmp_794 = and_1766_cse | nor_tmp_137;
  assign mux_tmp_755 = MUX_s_1_2_2(or_tmp_794, or_tmp_793, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign mux_759_nl = MUX_s_1_2_2(mux_tmp_755, mux_tmp_754, or_tmp_731);
  assign or_1246_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_757 = MUX_s_1_2_2(mux_759_nl, or_1246_nl, ac_float_cctor_operator_return_sva);
  assign or_1251_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | mux_tmp_757;
  assign mux_tmp_758 = MUX_s_1_2_2(mux_tmp_757, or_1251_nl, and_dcpl_1295);
  assign or_1252_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_758;
  assign mux_tmp_759 = MUX_s_1_2_2(mux_tmp_758, or_1252_nl, and_dcpl_1332);
  assign or_1253_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | mux_tmp_759;
  assign mux_tmp_760 = MUX_s_1_2_2(mux_tmp_759, or_1253_nl, and_dcpl_1304);
  assign or_1254_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_760;
  assign mux_tmp_761 = MUX_s_1_2_2(mux_tmp_760, or_1254_nl, and_dcpl_1291);
  assign or_1255_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | mux_tmp_761;
  assign mux_tmp_762 = MUX_s_1_2_2(mux_tmp_761, or_1255_nl, and_dcpl_1307);
  assign or_1256_nl = or_tmp_783 | mux_tmp_762;
  assign mux_tmp_763 = MUX_s_1_2_2(mux_tmp_762, or_1256_nl, and_dcpl_101);
  assign or_1257_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_763;
  assign mux_tmp_764 = MUX_s_1_2_2(mux_tmp_763, or_1257_nl, and_dcpl_1287);
  assign or_1258_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_operator_return_9_sva | mux_tmp_764;
  assign mux_tmp_765 = MUX_s_1_2_2(mux_tmp_764, or_1258_nl, and_dcpl_1298);
  assign or_1259_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_765;
  assign mux_tmp_766 = MUX_s_1_2_2(mux_tmp_765, or_1259_nl, and_dcpl_1338);
  assign or_1260_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_766;
  assign mux_tmp_767 = MUX_s_1_2_2(mux_tmp_766, or_1260_nl, and_dcpl_1344);
  assign or_1262_nl = and_dcpl_108 | mux_tmp_732;
  assign or_1261_nl = and_dcpl_108 | mux_tmp_767;
  assign mux_tmp_768 = MUX_s_1_2_2(or_1262_nl, or_1261_nl, and_dcpl_919);
  assign mux_772_nl = MUX_s_1_2_2(mux_tmp_768, or_tmp_747, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1263_nl = or_tmp_748 | mux_772_nl;
  assign mux_tmp_770 = MUX_s_1_2_2(mux_tmp_768, or_1263_nl, and_dcpl_1335);
  assign mux_tmp_771 = MUX_s_1_2_2(mux_tmp_770, mux_tmp_733, or_tmp_777);
  assign mux_tmp_772 = MUX_s_1_2_2(mux_tmp_752, mux_tmp_733, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_773 = MUX_s_1_2_2(or_tmp_792, or_tmp_734, or_tmp_762);
  assign mux_tmp_774 = MUX_s_1_2_2(or_tmp_792, or_tmp_734, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm);
  assign mux_tmp_775 = MUX_s_1_2_2(or_tmp_794, or_tmp_793, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm);
  assign mux_tmp_776 = MUX_s_1_2_2(mux_tmp_775, mux_tmp_774, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva);
  assign or_1281_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_777 = MUX_s_1_2_2(mux_tmp_776, or_1281_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign mux_781_nl = MUX_s_1_2_2(mux_tmp_777, mux_tmp_773, or_tmp_731);
  assign or_1277_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_779 = MUX_s_1_2_2(mux_781_nl, or_1277_nl, ac_float_cctor_operator_return_sva);
  assign or_1282_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_779;
  assign mux_tmp_780 = MUX_s_1_2_2(mux_tmp_779, or_1282_nl, and_dcpl_1295);
  assign or_1283_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_780;
  assign mux_tmp_781 = MUX_s_1_2_2(mux_tmp_780, or_1283_nl, and_dcpl_1332);
  assign or_1284_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_781;
  assign mux_tmp_782 = MUX_s_1_2_2(mux_tmp_781, or_1284_nl, and_dcpl_1304);
  assign or_1285_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_782;
  assign mux_tmp_783 = MUX_s_1_2_2(mux_tmp_782, or_1285_nl, and_dcpl_1291);
  assign or_1286_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_783;
  assign mux_tmp_784 = MUX_s_1_2_2(mux_tmp_783, or_1286_nl, and_dcpl_1307);
  assign or_1287_nl = or_tmp_783 | mux_tmp_784;
  assign mux_tmp_785 = MUX_s_1_2_2(mux_tmp_784, or_1287_nl, and_dcpl_101);
  assign or_1288_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_785;
  assign mux_tmp_786 = MUX_s_1_2_2(mux_tmp_785, or_1288_nl, and_dcpl_1287);
  assign or_1289_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_operator_return_9_sva | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_786;
  assign mux_tmp_787 = MUX_s_1_2_2(mux_tmp_786, or_1289_nl, and_dcpl_1298);
  assign or_1290_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_787;
  assign mux_tmp_788 = MUX_s_1_2_2(mux_tmp_787, or_1290_nl, and_dcpl_1338);
  assign or_1291_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_788;
  assign mux_792_nl = MUX_s_1_2_2(mux_tmp_788, or_1291_nl, and_dcpl_1344);
  assign mux_793_nl = MUX_s_1_2_2(mux_tmp_767, mux_792_nl, and_dcpl_108);
  assign mux_tmp_791 = MUX_s_1_2_2(mux_tmp_750, mux_793_nl, and_dcpl_919);
  assign mux_795_nl = MUX_s_1_2_2(mux_tmp_791, mux_tmp_768, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign mux_796_nl = MUX_s_1_2_2(mux_795_nl, mux_tmp_751, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1292_nl = or_tmp_748 | mux_796_nl;
  assign mux_tmp_794 = MUX_s_1_2_2(mux_tmp_791, or_1292_nl, and_dcpl_1335);
  assign mux_tmp_795 = MUX_s_1_2_2(mux_tmp_794, mux_tmp_770, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_796 = MUX_s_1_2_2(mux_tmp_795, mux_tmp_772, or_tmp_777);
  assign or_tmp_838 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm;
  assign mux_tmp_801 = MUX_s_1_2_2(mux_tmp_795, mux_tmp_772, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_tmp_809 = MUX_s_1_2_2(mux_tmp_770, mux_tmp_733, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign mux_tmp_810 = MUX_s_1_2_2(mux_tmp_794, mux_tmp_752, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign and_1781_cse = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      & and_dcpl_1301;
  assign and_1775_cse = and_dcpl_101 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva;
  assign or_1309_nl = and_1781_cse | and_dcpl_1347;
  assign mux_824_nl = MUX_s_1_2_2(and_1781_cse, or_1309_nl, ac_float_cctor_operator_return_sva);
  assign or_tmp_863 = (and_dcpl_1344 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm)
      | (and_dcpl_1338 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm)
      | (and_dcpl_1298 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva)
      | (and_dcpl_1287 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva)
      | and_1775_cse | (and_dcpl_1307 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva)
      | (and_dcpl_1291 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva)
      | (and_dcpl_1304 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva)
      | (and_dcpl_1332 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm)
      | (and_dcpl_1295 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva)
      | mux_824_nl;
  assign or_tmp_864 = (and_dcpl_1335 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm)
      | and_dcpl_919 | and_dcpl_108 | or_tmp_863;
  assign or_tmp_866 = or_tmp_746 | or_tmp_863;
  assign or_tmp_876 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva;
  assign mux_825_nl = MUX_s_1_2_2(nor_tmp_135, mux_tmp_735, or_tmp_876);
  assign or_1333_nl = (or_tmp_876 & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_823 = MUX_s_1_2_2(mux_825_nl, or_1333_nl, ac_float_cctor_operator_return_sva);
  assign or_1335_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_823;
  assign mux_tmp_824 = MUX_s_1_2_2(mux_tmp_823, or_1335_nl, and_dcpl_1295);
  assign or_1336_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_824;
  assign mux_tmp_825 = MUX_s_1_2_2(mux_tmp_824, or_1336_nl, and_dcpl_1332);
  assign or_1337_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_825;
  assign mux_tmp_826 = MUX_s_1_2_2(mux_tmp_825, or_1337_nl, and_dcpl_1304);
  assign or_1338_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | mux_tmp_826;
  assign mux_tmp_827 = MUX_s_1_2_2(mux_tmp_826, or_1338_nl, and_dcpl_1291);
  assign or_1339_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_827;
  assign mux_831_nl = MUX_s_1_2_2(mux_tmp_827, or_1339_nl, and_dcpl_1307);
  assign or_tmp_884 = and_1775_cse | mux_831_nl;
  assign or_1341_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | or_tmp_884;
  assign mux_tmp_829 = MUX_s_1_2_2(or_tmp_884, or_1341_nl, and_dcpl_1287);
  assign or_1342_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_829;
  assign mux_tmp_830 = MUX_s_1_2_2(mux_tmp_829, or_1342_nl, and_dcpl_1298);
  assign or_1343_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_830;
  assign mux_tmp_831 = MUX_s_1_2_2(mux_tmp_830, or_1343_nl, and_dcpl_1338);
  assign or_1344_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | mux_tmp_831;
  assign mux_835_nl = MUX_s_1_2_2(mux_tmp_831, or_1344_nl, and_dcpl_1344);
  assign mux_tmp_833 = MUX_s_1_2_2(or_tmp_863, mux_835_nl, and_dcpl_108);
  assign or_tmp_889 = and_dcpl_919 | mux_tmp_833;
  assign mux_tmp_834 = MUX_s_1_2_2(or_tmp_889, or_tmp_866, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign or_1346_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | mux_tmp_834;
  assign mux_tmp_835 = MUX_s_1_2_2(or_tmp_889, or_1346_nl, and_dcpl_1335);
  assign or_tmp_897 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva;
  assign and_1786_cse = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      & and_dcpl_1301;
  assign or_1362_nl = and_1786_cse | nor_tmp_137;
  assign or_1360_nl = and_1786_cse | and_dcpl_1347;
  assign mux_tmp_837 = MUX_s_1_2_2(or_1362_nl, or_1360_nl, ac_float_cctor_operator_return_sva);
  assign or_1363_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | mux_tmp_837;
  assign mux_tmp_838 = MUX_s_1_2_2(mux_tmp_837, or_1363_nl, and_dcpl_1295);
  assign or_1364_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_838;
  assign mux_tmp_839 = MUX_s_1_2_2(mux_tmp_838, or_1364_nl, and_dcpl_1332);
  assign or_1365_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | mux_tmp_839;
  assign mux_tmp_840 = MUX_s_1_2_2(mux_tmp_839, or_1365_nl, and_dcpl_1304);
  assign or_1366_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_840;
  assign mux_tmp_841 = MUX_s_1_2_2(mux_tmp_840, or_1366_nl, and_dcpl_1291);
  assign or_1367_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | mux_tmp_841;
  assign mux_tmp_842 = MUX_s_1_2_2(mux_tmp_841, or_1367_nl, and_dcpl_1307);
  assign or_1368_nl = or_tmp_897 | mux_tmp_842;
  assign mux_tmp_843 = MUX_s_1_2_2(mux_tmp_842, or_1368_nl, and_dcpl_101);
  assign or_1369_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | mux_tmp_843;
  assign mux_tmp_844 = MUX_s_1_2_2(mux_tmp_843, or_1369_nl, and_dcpl_1287);
  assign or_1370_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_operator_return_9_sva | mux_tmp_844;
  assign mux_tmp_845 = MUX_s_1_2_2(mux_tmp_844, or_1370_nl, and_dcpl_1298);
  assign or_1371_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_845;
  assign mux_tmp_846 = MUX_s_1_2_2(mux_tmp_845, or_1371_nl, and_dcpl_1338);
  assign or_1372_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_846;
  assign mux_tmp_847 = MUX_s_1_2_2(mux_tmp_846, or_1372_nl, and_dcpl_1344);
  assign or_1374_nl = and_dcpl_108 | or_tmp_863;
  assign or_1373_nl = and_dcpl_108 | mux_tmp_847;
  assign mux_tmp_848 = MUX_s_1_2_2(or_1374_nl, or_1373_nl, and_dcpl_919);
  assign mux_852_nl = MUX_s_1_2_2(mux_tmp_848, or_tmp_866, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1375_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | mux_852_nl;
  assign mux_tmp_850 = MUX_s_1_2_2(mux_tmp_848, or_1375_nl, and_dcpl_1335);
  assign mux_tmp_851 = MUX_s_1_2_2(mux_tmp_850, or_tmp_864, or_tmp_777);
  assign mux_tmp_852 = MUX_s_1_2_2(mux_tmp_835, or_tmp_864, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_856_nl = MUX_s_1_2_2(mux_tmp_775, mux_tmp_774, or_tmp_876);
  assign or_1388_nl = ((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva)
      & and_dcpl_1301) | and_dcpl_1347;
  assign mux_tmp_854 = MUX_s_1_2_2(mux_856_nl, or_1388_nl, ac_float_cctor_operator_return_sva);
  assign or_1390_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_854;
  assign mux_tmp_855 = MUX_s_1_2_2(mux_tmp_854, or_1390_nl, and_dcpl_1295);
  assign or_1391_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | mux_tmp_855;
  assign mux_tmp_856 = MUX_s_1_2_2(mux_tmp_855, or_1391_nl, and_dcpl_1332);
  assign or_1392_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_856;
  assign mux_tmp_857 = MUX_s_1_2_2(mux_tmp_856, or_1392_nl, and_dcpl_1304);
  assign or_1393_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_857;
  assign mux_tmp_858 = MUX_s_1_2_2(mux_tmp_857, or_1393_nl, and_dcpl_1291);
  assign or_1394_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_858;
  assign mux_tmp_859 = MUX_s_1_2_2(mux_tmp_858, or_1394_nl, and_dcpl_1307);
  assign or_1395_nl = or_tmp_897 | mux_tmp_859;
  assign mux_tmp_860 = MUX_s_1_2_2(mux_tmp_859, or_1395_nl, and_dcpl_101);
  assign or_1396_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | mux_tmp_860;
  assign mux_tmp_861 = MUX_s_1_2_2(mux_tmp_860, or_1396_nl, and_dcpl_1287);
  assign or_1397_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | ac_float_cctor_operator_return_9_sva | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_861;
  assign mux_tmp_862 = MUX_s_1_2_2(mux_tmp_861, or_1397_nl, and_dcpl_1298);
  assign or_1398_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
      | mux_tmp_862;
  assign mux_tmp_863 = MUX_s_1_2_2(mux_tmp_862, or_1398_nl, and_dcpl_1338);
  assign or_1399_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_863;
  assign mux_867_nl = MUX_s_1_2_2(mux_tmp_863, or_1399_nl, and_dcpl_1344);
  assign mux_868_nl = MUX_s_1_2_2(mux_tmp_847, mux_867_nl, and_dcpl_108);
  assign mux_tmp_866 = MUX_s_1_2_2(mux_tmp_833, mux_868_nl, and_dcpl_919);
  assign mux_870_nl = MUX_s_1_2_2(mux_tmp_866, mux_tmp_848, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign mux_871_nl = MUX_s_1_2_2(mux_870_nl, mux_tmp_834, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1400_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | mux_871_nl;
  assign mux_tmp_869 = MUX_s_1_2_2(mux_tmp_866, or_1400_nl, and_dcpl_1335);
  assign mux_tmp_870 = MUX_s_1_2_2(mux_tmp_869, mux_tmp_850, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_871 = MUX_s_1_2_2(mux_tmp_870, mux_tmp_852, or_tmp_777);
  assign mux_tmp_876 = MUX_s_1_2_2(mux_tmp_870, mux_tmp_852, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_tmp_884 = MUX_s_1_2_2(mux_tmp_850, or_tmp_864, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign mux_tmp_885 = MUX_s_1_2_2(mux_tmp_869, mux_tmp_835, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign and_1793_cse = and_dcpl_101 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  assign mux_904_nl = MUX_s_1_2_2(nor_tmp_132, mux_tmp, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva);
  assign or_tmp_970 = (and_dcpl_1344 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm)
      | (and_dcpl_1338 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm)
      | (and_dcpl_1298 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva)
      | (and_dcpl_1287 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva)
      | and_1793_cse | (and_dcpl_1307 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva)
      | (and_dcpl_1291 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva)
      | (and_dcpl_1304 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva)
      | (and_dcpl_1332 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm)
      | (and_dcpl_1295 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva)
      | mux_904_nl;
  assign or_tmp_971 = (and_dcpl_1335 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm)
      | and_dcpl_919 | and_dcpl_108 | or_tmp_970;
  assign or_tmp_973 = or_tmp_746 | or_tmp_970;
  assign mux_tmp_902 = MUX_s_1_2_2(mux_tmp_737, mux_tmp_734, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva);
  assign or_1439_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_902;
  assign mux_tmp_903 = MUX_s_1_2_2(mux_tmp_902, or_1439_nl, and_dcpl_1295);
  assign or_1440_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | mux_tmp_903;
  assign mux_tmp_904 = MUX_s_1_2_2(mux_tmp_903, or_1440_nl, and_dcpl_1332);
  assign or_1441_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_904;
  assign mux_tmp_905 = MUX_s_1_2_2(mux_tmp_904, or_1441_nl, and_dcpl_1304);
  assign or_1442_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | mux_tmp_905;
  assign mux_tmp_906 = MUX_s_1_2_2(mux_tmp_905, or_1442_nl, and_dcpl_1291);
  assign or_1443_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_906;
  assign mux_910_nl = MUX_s_1_2_2(mux_tmp_906, or_1443_nl, and_dcpl_1307);
  assign or_tmp_988 = and_1793_cse | mux_910_nl;
  assign or_1445_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | or_tmp_988;
  assign mux_tmp_908 = MUX_s_1_2_2(or_tmp_988, or_1445_nl, and_dcpl_1287);
  assign or_1446_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_908;
  assign mux_tmp_909 = MUX_s_1_2_2(mux_tmp_908, or_1446_nl, and_dcpl_1298);
  assign or_1447_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | mux_tmp_909;
  assign mux_tmp_910 = MUX_s_1_2_2(mux_tmp_909, or_1447_nl, and_dcpl_1338);
  assign or_1448_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | mux_tmp_910;
  assign mux_914_nl = MUX_s_1_2_2(mux_tmp_910, or_1448_nl, and_dcpl_1344);
  assign mux_tmp_912 = MUX_s_1_2_2(or_tmp_970, mux_914_nl, and_dcpl_108);
  assign or_tmp_993 = and_dcpl_919 | mux_tmp_912;
  assign mux_tmp_913 = MUX_s_1_2_2(or_tmp_993, or_tmp_973, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign or_1450_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
      | mux_tmp_913;
  assign mux_tmp_914 = MUX_s_1_2_2(or_tmp_993, or_1450_nl, and_dcpl_1335);
  assign or_tmp_1001 = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva;
  assign mux_tmp_916 = MUX_s_1_2_2(mux_tmp_755, mux_tmp_754, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva);
  assign or_1463_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | mux_tmp_916;
  assign mux_tmp_917 = MUX_s_1_2_2(mux_tmp_916, or_1463_nl, and_dcpl_1295);
  assign or_1464_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | mux_tmp_917;
  assign mux_tmp_918 = MUX_s_1_2_2(mux_tmp_917, or_1464_nl, and_dcpl_1332);
  assign or_1465_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | mux_tmp_918;
  assign mux_tmp_919 = MUX_s_1_2_2(mux_tmp_918, or_1465_nl, and_dcpl_1304);
  assign or_1466_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_919;
  assign mux_tmp_920 = MUX_s_1_2_2(mux_tmp_919, or_1466_nl, and_dcpl_1291);
  assign or_1467_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | mux_tmp_920;
  assign mux_tmp_921 = MUX_s_1_2_2(mux_tmp_920, or_1467_nl, and_dcpl_1307);
  assign or_1468_nl = or_tmp_1001 | mux_tmp_921;
  assign mux_tmp_922 = MUX_s_1_2_2(mux_tmp_921, or_1468_nl, and_dcpl_101);
  assign or_1469_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_922;
  assign mux_tmp_923 = MUX_s_1_2_2(mux_tmp_922, or_1469_nl, and_dcpl_1287);
  assign or_1470_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_operator_return_9_sva | mux_tmp_923;
  assign mux_tmp_924 = MUX_s_1_2_2(mux_tmp_923, or_1470_nl, and_dcpl_1298);
  assign or_1471_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | mux_tmp_924;
  assign mux_tmp_925 = MUX_s_1_2_2(mux_tmp_924, or_1471_nl, and_dcpl_1338);
  assign or_1472_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_925;
  assign mux_tmp_926 = MUX_s_1_2_2(mux_tmp_925, or_1472_nl, and_dcpl_1344);
  assign or_1474_nl = and_dcpl_108 | or_tmp_970;
  assign or_1473_nl = and_dcpl_108 | mux_tmp_926;
  assign mux_tmp_927 = MUX_s_1_2_2(or_1474_nl, or_1473_nl, and_dcpl_919);
  assign mux_931_nl = MUX_s_1_2_2(mux_tmp_927, or_tmp_973, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1475_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
      | mux_931_nl;
  assign mux_tmp_929 = MUX_s_1_2_2(mux_tmp_927, or_1475_nl, and_dcpl_1335);
  assign mux_tmp_930 = MUX_s_1_2_2(mux_tmp_929, or_tmp_971, or_tmp_777);
  assign mux_tmp_931 = MUX_s_1_2_2(mux_tmp_914, or_tmp_971, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_932 = MUX_s_1_2_2(mux_tmp_777, mux_tmp_773, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva);
  assign or_1487_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_932;
  assign mux_tmp_933 = MUX_s_1_2_2(mux_tmp_932, or_1487_nl, and_dcpl_1295);
  assign or_1488_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | mux_tmp_933;
  assign mux_tmp_934 = MUX_s_1_2_2(mux_tmp_933, or_1488_nl, and_dcpl_1332);
  assign or_1489_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_934;
  assign mux_tmp_935 = MUX_s_1_2_2(mux_tmp_934, or_1489_nl, and_dcpl_1304);
  assign or_1490_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_935;
  assign mux_tmp_936 = MUX_s_1_2_2(mux_tmp_935, or_1490_nl, and_dcpl_1291);
  assign or_1491_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_936;
  assign mux_tmp_937 = MUX_s_1_2_2(mux_tmp_936, or_1491_nl, and_dcpl_1307);
  assign or_1492_nl = or_tmp_1001 | mux_tmp_937;
  assign mux_tmp_938 = MUX_s_1_2_2(mux_tmp_937, or_1492_nl, and_dcpl_101);
  assign or_1493_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | mux_tmp_938;
  assign mux_tmp_939 = MUX_s_1_2_2(mux_tmp_938, or_1493_nl, and_dcpl_1287);
  assign or_1494_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | ac_float_cctor_operator_return_9_sva | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_939;
  assign mux_tmp_940 = MUX_s_1_2_2(mux_tmp_939, or_1494_nl, and_dcpl_1298);
  assign or_1495_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
      | mux_tmp_940;
  assign mux_tmp_941 = MUX_s_1_2_2(mux_tmp_940, or_1495_nl, and_dcpl_1338);
  assign or_1496_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_941;
  assign mux_945_nl = MUX_s_1_2_2(mux_tmp_941, or_1496_nl, and_dcpl_1344);
  assign mux_946_nl = MUX_s_1_2_2(mux_tmp_926, mux_945_nl, and_dcpl_108);
  assign mux_tmp_944 = MUX_s_1_2_2(mux_tmp_912, mux_946_nl, and_dcpl_919);
  assign mux_948_nl = MUX_s_1_2_2(mux_tmp_944, mux_tmp_927, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign mux_949_nl = MUX_s_1_2_2(mux_948_nl, mux_tmp_913, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign or_1497_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
      | mux_949_nl;
  assign mux_tmp_947 = MUX_s_1_2_2(mux_tmp_944, or_1497_nl, and_dcpl_1335);
  assign mux_tmp_948 = MUX_s_1_2_2(mux_tmp_947, mux_tmp_929, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_949 = MUX_s_1_2_2(mux_tmp_948, mux_tmp_931, or_tmp_777);
  assign mux_tmp_954 = MUX_s_1_2_2(mux_tmp_948, mux_tmp_931, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_tmp_962 = MUX_s_1_2_2(mux_tmp_929, or_tmp_971, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign mux_tmp_963 = MUX_s_1_2_2(mux_tmp_947, mux_tmp_914, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign and_tmp_29 = and_dcpl_108 & ((and_dcpl_1344 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm)
      | (and_dcpl_1338 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm)
      | (and_dcpl_1298 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva)
      | (and_dcpl_1287 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva)
      | (and_dcpl_1307 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva)
      | (and_dcpl_1291 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm)
      | (and_dcpl_1304 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva)
      | (and_dcpl_1332 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva)
      | (and_dcpl_1295 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm)
      | mux_tmp_736);
  assign or_tmp_1062 = and_dcpl_919 | and_tmp_29;
  assign and_1815_cse = and_dcpl_101 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva;
  assign or_tmp_1074 = (and_dcpl_1344 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm)
      | (and_dcpl_1338 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm)
      | (and_dcpl_1298 & ac_float_cctor_operator_return_9_sva) | (and_dcpl_1287 &
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva)
      | and_1815_cse | (and_dcpl_1307 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva)
      | (and_dcpl_1291 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm)
      | (and_dcpl_1304 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva)
      | (and_dcpl_1332 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva)
      | (and_dcpl_1295 & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm)
      | or_tmp_794;
  assign or_1531_nl = and_dcpl_108 | or_tmp_1074;
  assign mux_tmp_976 = MUX_s_1_2_2(and_dcpl_108, or_1531_nl, and_dcpl_919);
  assign mux_1112_nl = MUX_s_1_2_2(mux_tmp_976, or_tmp_746, and_1829_cse);
  assign mux_tmp_978 = MUX_s_1_2_2(mux_1112_nl, or_tmp_746, or_tmp_777);
  assign mux_1117_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_tmp_979 = MUX_s_1_2_2(mux_1117_nl, or_tmp_746, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign or_1542_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | mux_tmp_776;
  assign mux_tmp_981 = MUX_s_1_2_2(mux_tmp_776, or_1542_nl, and_dcpl_1295);
  assign or_1543_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
      | mux_tmp_981;
  assign mux_tmp_982 = MUX_s_1_2_2(mux_tmp_981, or_1543_nl, and_dcpl_1332);
  assign or_1544_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | mux_tmp_982;
  assign mux_tmp_983 = MUX_s_1_2_2(mux_tmp_982, or_1544_nl, and_dcpl_1304);
  assign or_1545_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | mux_tmp_983;
  assign mux_tmp_984 = MUX_s_1_2_2(mux_tmp_983, or_1545_nl, and_dcpl_1291);
  assign or_1546_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | mux_tmp_984;
  assign mux_988_nl = MUX_s_1_2_2(mux_tmp_984, or_1546_nl, and_dcpl_1307);
  assign or_tmp_1091 = and_1815_cse | mux_988_nl;
  assign or_1548_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | or_tmp_1091;
  assign mux_tmp_986 = MUX_s_1_2_2(or_tmp_1091, or_1548_nl, and_dcpl_1287);
  assign or_1549_nl = ac_float_cctor_operator_return_9_sva | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | mux_tmp_986;
  assign mux_tmp_987 = MUX_s_1_2_2(mux_tmp_986, or_1549_nl, and_dcpl_1298);
  assign or_1550_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | mux_tmp_987;
  assign mux_tmp_988 = MUX_s_1_2_2(mux_tmp_987, or_1550_nl, and_dcpl_1338);
  assign or_1551_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | mux_tmp_988;
  assign mux_992_nl = MUX_s_1_2_2(mux_tmp_988, or_1551_nl, and_dcpl_1344);
  assign mux_993_nl = MUX_s_1_2_2(or_tmp_1074, mux_992_nl, and_dcpl_108);
  assign mux_tmp_991 = MUX_s_1_2_2(and_tmp_29, mux_993_nl, and_dcpl_919);
  assign mux_995_nl = MUX_s_1_2_2(mux_tmp_991, mux_tmp_976, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign mux_983_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign mux_996_nl = MUX_s_1_2_2(mux_995_nl, mux_983_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm);
  assign mux_tmp_994 = MUX_s_1_2_2(mux_tmp_991, mux_996_nl, and_dcpl_1335);
  assign mux_tmp_995 = MUX_s_1_2_2(mux_tmp_994, mux_1035_itm, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm);
  assign mux_tmp_996 = MUX_s_1_2_2(mux_tmp_995, mux_tmp_979, or_tmp_777);
  assign mux_tmp_1001 = MUX_s_1_2_2(mux_tmp_995, mux_tmp_979, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm);
  assign mux_1113_nl = MUX_s_1_2_2(mux_tmp_976, or_tmp_746, and_1829_cse);
  assign mux_tmp_1009 = MUX_s_1_2_2(mux_1113_nl, or_tmp_746, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign mux_1039_nl = MUX_s_1_2_2(or_tmp_1062, or_tmp_746, and_1827_cse);
  assign mux_tmp_1010 = MUX_s_1_2_2(mux_tmp_994, mux_1039_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign nor_773_cse = ~((fsm_output[7]) | (fsm_output[3]) | (fsm_output[5]));
  assign nor_774_cse = ~((fsm_output[4]) | (fsm_output[8]));
  assign and_dcpl_1635 = nor_773_cse & nor_774_cse;
  assign and_dcpl_1640 = and_dcpl_1635 & nor_221_cse & (fsm_output[2]) & (~ (fsm_output[6]));
  assign and_dcpl_1663 = nor_773_cse & nor_774_cse & nor_221_cse & (fsm_output[2])
      & (~ (fsm_output[6]));
  assign and_568_ssc = and_dcpl_102 & ((operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1!=2'b00))
      & (~((fsm_output[0]) | (fsm_output[6]))) & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp
      & (~ operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0) & (fsm_output[3:2]==2'b01)
      & and_dcpl_85;
  assign and_573_ssc = (MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_cse
      | (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp) | operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0)
      & and_dcpl_103 & and_dcpl_547;
  assign or_242_nl = (fsm_output[1:0]!=2'b01);
  assign mux_318_nl = MUX_s_1_2_2(or_242_nl, mux_tmp_314, nor_68_cse);
  assign mux_319_nl = MUX_s_1_2_2(mux_318_nl, mux_tmp_314, MAC_3_result_operator_result_operator_nor_tmp);
  assign and_575_ssc = (~(mux_319_nl | (fsm_output[8]))) & and_dcpl_547;
  assign mux_390_nl = MUX_s_1_2_2(nor_369_cse, (fsm_output[7]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva);
  assign or_563_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      | (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_562_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
      | (~ (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_389_nl = MUX_s_1_2_2(or_563_nl, or_562_nl, fsm_output[7]);
  assign mux_391_nl = MUX_s_1_2_2(mux_390_nl, mux_389_nl, fsm_output[5]);
  assign nor_371_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
      | (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_386_nl = MUX_s_1_2_2(or_tmp_374, nor_371_nl, MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_387_nl = MUX_s_1_2_2(mux_386_nl, or_tmp_374, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva);
  assign nor_373_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
      | (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_384_nl = MUX_s_1_2_2(or_tmp_370, nor_373_nl, MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_385_nl = MUX_s_1_2_2(mux_384_nl, or_tmp_370, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm);
  assign mux_388_nl = MUX_s_1_2_2(mux_387_nl, mux_385_nl, fsm_output[5]);
  assign mux_392_nl = MUX_s_1_2_2(mux_391_nl, mux_388_nl, fsm_output[4]);
  assign or_553_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
      | (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_552_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
      | (~ (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_381_nl = MUX_s_1_2_2(or_553_nl, or_552_nl, fsm_output[7]);
  assign or_551_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
      | (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_550_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
      | (~ (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_380_nl = MUX_s_1_2_2(or_551_nl, or_550_nl, fsm_output[7]);
  assign mux_382_nl = MUX_s_1_2_2(mux_381_nl, mux_380_nl, fsm_output[5]);
  assign nor_375_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
      | (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_377_nl = MUX_s_1_2_2(or_tmp_362, nor_375_nl, MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_378_nl = MUX_s_1_2_2(mux_377_nl, or_tmp_362, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm);
  assign or_545_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
      | (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_544_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm
      | (~ (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_376_nl = MUX_s_1_2_2(or_545_nl, or_544_nl, fsm_output[7]);
  assign mux_379_nl = MUX_s_1_2_2(mux_378_nl, mux_376_nl, fsm_output[5]);
  assign mux_383_nl = MUX_s_1_2_2(mux_382_nl, mux_379_nl, fsm_output[4]);
  assign mux_393_nl = MUX_s_1_2_2(mux_392_nl, mux_383_nl, fsm_output[3]);
  assign nor_377_nl = ~((fsm_output[7]) | nor_68_cse);
  assign mux_371_nl = MUX_s_1_2_2(or_tmp_356, nor_377_nl, MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_372_nl = MUX_s_1_2_2(mux_371_nl, or_tmp_356, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva);
  assign or_539_nl = ac_float_cctor_operator_return_9_sva | (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_538_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
      | (~ (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_370_nl = MUX_s_1_2_2(or_539_nl, or_538_nl, fsm_output[7]);
  assign mux_373_nl = MUX_s_1_2_2(mux_372_nl, mux_370_nl, fsm_output[5]);
  assign or_537_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
      | (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_536_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
      | (~ (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_368_nl = MUX_s_1_2_2(or_537_nl, or_536_nl, fsm_output[7]);
  assign or_535_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
      | (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_534_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
      | (~ (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_367_nl = MUX_s_1_2_2(or_535_nl, or_534_nl, fsm_output[7]);
  assign mux_369_nl = MUX_s_1_2_2(mux_368_nl, mux_367_nl, fsm_output[5]);
  assign mux_374_nl = MUX_s_1_2_2(mux_373_nl, mux_369_nl, fsm_output[4]);
  assign nor_379_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
      | (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_363_nl = MUX_s_1_2_2(or_tmp_346, nor_379_nl, MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_364_nl = MUX_s_1_2_2(mux_363_nl, or_tmp_346, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva);
  assign or_529_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
      | (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_528_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm
      | (~ (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_362_nl = MUX_s_1_2_2(or_529_nl, or_528_nl, fsm_output[7]);
  assign mux_365_nl = MUX_s_1_2_2(mux_364_nl, mux_362_nl, fsm_output[5]);
  assign or_527_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
      | (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_526_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
      | (~ (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_360_nl = MUX_s_1_2_2(or_527_nl, or_526_nl, fsm_output[7]);
  assign or_525_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
      | (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_524_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm
      | (~ (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_359_nl = MUX_s_1_2_2(or_525_nl, or_524_nl, fsm_output[7]);
  assign mux_361_nl = MUX_s_1_2_2(mux_360_nl, mux_359_nl, fsm_output[5]);
  assign mux_366_nl = MUX_s_1_2_2(mux_365_nl, mux_361_nl, fsm_output[4]);
  assign mux_375_nl = MUX_s_1_2_2(mux_374_nl, mux_366_nl, fsm_output[3]);
  assign mux_394_nl = MUX_s_1_2_2(mux_393_nl, mux_375_nl, fsm_output[2]);
  assign or_523_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva
      | (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_522_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
      | (~ (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_354_nl = MUX_s_1_2_2(or_523_nl, or_522_nl, fsm_output[7]);
  assign nor_381_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
      | (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_352_nl = MUX_s_1_2_2(or_tmp_334, nor_381_nl, MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_353_nl = MUX_s_1_2_2(mux_352_nl, or_tmp_334, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm);
  assign mux_355_nl = MUX_s_1_2_2(mux_354_nl, mux_353_nl, fsm_output[5]);
  assign nor_383_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
      | (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_349_nl = MUX_s_1_2_2(or_tmp_330, nor_383_nl, MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_350_nl = MUX_s_1_2_2(mux_349_nl, or_tmp_330, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm);
  assign nor_385_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
      | (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_347_nl = MUX_s_1_2_2(or_tmp_326, nor_385_nl, MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_348_nl = MUX_s_1_2_2(mux_347_nl, or_tmp_326, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign mux_351_nl = MUX_s_1_2_2(mux_350_nl, mux_348_nl, fsm_output[5]);
  assign mux_356_nl = MUX_s_1_2_2(mux_355_nl, mux_351_nl, fsm_output[4]);
  assign or_509_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_508_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
      | (~ (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_344_nl = MUX_s_1_2_2(or_509_nl, or_508_nl, fsm_output[7]);
  assign or_507_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
      | (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_506_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm
      | (~ (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_343_nl = MUX_s_1_2_2(or_507_nl, or_506_nl, fsm_output[7]);
  assign mux_345_nl = MUX_s_1_2_2(mux_344_nl, mux_343_nl, fsm_output[5]);
  assign nor_387_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
      | (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_340_nl = MUX_s_1_2_2(or_tmp_318, nor_387_nl, MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_341_nl = MUX_s_1_2_2(mux_340_nl, or_tmp_318, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm);
  assign nor_389_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
      | (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_338_nl = MUX_s_1_2_2(or_tmp_314, nor_389_nl, MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_339_nl = MUX_s_1_2_2(mux_338_nl, or_tmp_314, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign mux_342_nl = MUX_s_1_2_2(mux_341_nl, mux_339_nl, fsm_output[5]);
  assign mux_346_nl = MUX_s_1_2_2(mux_345_nl, mux_342_nl, fsm_output[4]);
  assign mux_357_nl = MUX_s_1_2_2(mux_356_nl, mux_346_nl, fsm_output[3]);
  assign or_497_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
      | (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_496_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
      | (~ (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_334_nl = MUX_s_1_2_2(or_497_nl, or_496_nl, fsm_output[7]);
  assign nor_391_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
      | (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_332_nl = MUX_s_1_2_2(or_tmp_308, nor_391_nl, MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_333_nl = MUX_s_1_2_2(mux_332_nl, or_tmp_308, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm);
  assign mux_335_nl = MUX_s_1_2_2(mux_334_nl, mux_333_nl, fsm_output[5]);
  assign or_491_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
      | (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_490_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
      | (~ (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_330_nl = MUX_s_1_2_2(or_491_nl, or_490_nl, fsm_output[7]);
  assign or_489_nl = (~ (fsm_output[7])) | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | (~ (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign and_578_nl = (fsm_output[7]) & (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
      | (~ (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign nor_70_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
      | (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])));
  assign mux_329_nl = MUX_s_1_2_2(or_489_nl, and_578_nl, nor_70_nl);
  assign mux_331_nl = MUX_s_1_2_2(mux_330_nl, mux_329_nl, fsm_output[5]);
  assign mux_336_nl = MUX_s_1_2_2(mux_335_nl, mux_331_nl, fsm_output[4]);
  assign or_486_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
      | (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_485_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm
      | (~ (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_326_nl = MUX_s_1_2_2(or_486_nl, or_485_nl, fsm_output[7]);
  assign nor_393_nl = ~((fsm_output[7]) | (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
      | (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])))));
  assign mux_324_nl = MUX_s_1_2_2(or_tmp_297, nor_393_nl, MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_325_nl = MUX_s_1_2_2(mux_324_nl, or_tmp_297, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign mux_327_nl = MUX_s_1_2_2(mux_326_nl, mux_325_nl, fsm_output[5]);
  assign or_480_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
      | (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign or_479_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | (~ (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]));
  assign mux_322_nl = MUX_s_1_2_2(or_480_nl, or_479_nl, fsm_output[7]);
  assign nor_394_nl = ~((~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
      | (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))))
      | (fsm_output[7]));
  assign mux_320_nl = MUX_s_1_2_2(or_tmp_292, nor_394_nl, MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]);
  assign mux_321_nl = MUX_s_1_2_2(mux_320_nl, or_tmp_292, ac_float_cctor_operator_return_sva);
  assign mux_323_nl = MUX_s_1_2_2(mux_322_nl, mux_321_nl, fsm_output[5]);
  assign mux_328_nl = MUX_s_1_2_2(mux_327_nl, mux_323_nl, fsm_output[4]);
  assign mux_337_nl = MUX_s_1_2_2(mux_336_nl, mux_328_nl, fsm_output[3]);
  assign mux_358_nl = MUX_s_1_2_2(mux_357_nl, mux_337_nl, fsm_output[2]);
  assign mux_395_nl = MUX_s_1_2_2(mux_394_nl, mux_358_nl, fsm_output[6]);
  assign and_579_ssc = mux_395_nl & and_dcpl_106 & (~((fsm_output[0]) | MAC_3_result_operator_result_operator_nor_tmp));
  assign and_584_ssc = (((MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_85;
  assign and_589_ssc = (((MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_85;
  assign and_595_ssc = (((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_567;
  assign and_599_ssc = (((MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_567;
  assign and_603_ssc = (((MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_567;
  assign and_607_ssc = (((MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_567;
  assign and_613_ssc = (((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_585;
  assign and_617_ssc = (((MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_9_sva)) | MAC_3_result_operator_result_operator_nor_tmp)
      & and_dcpl_107 & and_dcpl_546 & and_dcpl_585;
  assign and_621_ssc = (((MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_585;
  assign and_625_ssc = (((MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_585;
  assign and_631_ssc = (((MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_603;
  assign and_635_ssc = (((MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_603;
  assign and_639_ssc = (((MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_603;
  assign and_643_ssc = (((MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_603;
  assign and_649_ssc = (((MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_85;
  assign and_655_ssc = (((MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_85;
  assign and_660_ssc = (((MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_85;
  assign and_665_ssc = (((MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_85;
  assign and_669_ssc = (((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_567;
  assign and_673_ssc = (((MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_567;
  assign and_677_ssc = (((MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_567;
  assign and_681_ssc = (((MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_567;
  assign and_685_ssc = (((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_585;
  assign and_689_ssc = (((MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_585;
  assign and_693_ssc = (((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_585;
  assign and_697_ssc = (((MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_585;
  assign and_701_ssc = (((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_603;
  assign and_705_ssc = (((MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_603;
  assign and_709_ssc = (((MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_603;
  assign and_713_ssc = (((MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_603;
  assign and_718_ssc = (((MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_690;
  assign and_722_ssc = (((MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_690;
  assign and_726_ssc = (((MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_690;
  assign and_730_ssc = (((MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_690;
  assign and_735_ssc = (((MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_707;
  assign and_739_ssc = (((MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_707;
  assign and_743_ssc = (((MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_707;
  assign and_747_ssc = (((MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_707;
  assign and_752_ssc = (((MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_724;
  assign and_756_ssc = (((MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_724;
  assign and_760_ssc = (((MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_724;
  assign and_764_ssc = (((MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_724;
  assign and_769_ssc = (((MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_259
      & and_dcpl_741;
  assign and_773_ssc = (((MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_546
      & and_dcpl_741;
  assign and_777_ssc = (((MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_556
      & and_dcpl_741;
  assign and_781_ssc = (((MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_561
      & and_dcpl_741;
  assign and_785_ssc = (((MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_690;
  assign and_789_ssc = (((MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_690;
  assign and_793_ssc = (((MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_690;
  assign and_797_ssc = (((MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_690;
  assign and_801_ssc = (((MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_707;
  assign and_805_ssc = (((MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_707;
  assign and_809_ssc = (((MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_707;
  assign and_813_ssc = (((MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_707;
  assign and_817_ssc = (((MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_724;
  assign and_821_ssc = (((MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_724;
  assign and_825_ssc = (((MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_724;
  assign and_829_ssc = (((MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_637
      & and_dcpl_724;
  assign and_833_ssc = (((MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_621
      & and_dcpl_741;
  assign and_837_ssc = (((MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_627
      & and_dcpl_741;
  assign and_841_ssc = (((MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm))
      | MAC_3_result_operator_result_operator_nor_tmp) & and_dcpl_107 & and_dcpl_632
      & and_dcpl_741;
  assign and_845_ssc = (((MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & (~ ac_float_cctor_operator_return_sva)) | MAC_3_result_operator_result_operator_nor_tmp)
      & and_dcpl_107 & and_dcpl_637 & and_dcpl_741;
  assign nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt = conv_s2s_5_6(delay_lane_e_9_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[49:45]);
  assign MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt = nl_MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_95_itm
      = ~(and_dcpl_109 | ((or_dcpl_126 ^ (fsm_output[8])) & nor_221_cse));
  assign nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0 = conv_s2s_5_6(delay_lane_e_10_sva)
      + conv_s2s_5_6(taps_e_rsci_idat[54:50]);
  assign operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0 = nl_operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[5:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2}) + conv_s2s_6_7({1'b1
      , (~ MAC_1_leading_sign_18_1_1_0_cmp_rtn_oreg)}) + 7'b0000001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl[6:0];
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = ({operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1
      , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2}) + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_1_sva_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl
      = MUX_v_7_2_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_nl,
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva[21]))
      & MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl
      = MUX_v_7_2_2(7'b0000000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_nl);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0 + conv_u2s_4_7(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_2_sva_1);
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl
      = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl[6:0];
  assign and_1757_nl = and_dcpl_109 & (~ or_1557_tmp);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])))
      & and_dcpl_154;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_256_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1[1])
      & and_dcpl_154;
  assign operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0 = MUX1HOT_v_7_5_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl,
      z_out, MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_nl,
      7'b1110000, {and_dcpl_160 , and_1757_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_256_nl , or_1557_tmp});
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0
      = conv_s2s_5_6(delay_lane_e_40_sva) + conv_s2s_5_6(taps_e_rsci_idat[204:200]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0
      = conv_s2s_5_6(delay_lane_e_41_sva) + conv_s2s_5_6(taps_e_rsci_idat[209:205]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0
      = conv_s2s_5_6(delay_lane_e_42_sva) + conv_s2s_5_6(taps_e_rsci_idat[214:210]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0
      = conv_s2s_5_6(delay_lane_e_43_sva) + conv_s2s_5_6(taps_e_rsci_idat[219:215]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0
      = conv_s2s_5_6(delay_lane_e_44_sva) + conv_s2s_5_6(taps_e_rsci_idat[224:220]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0
      = conv_s2s_5_6(delay_lane_e_45_sva) + conv_s2s_5_6(taps_e_rsci_idat[229:225]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0
      = conv_s2s_5_6(delay_lane_e_46_sva) + conv_s2s_5_6(taps_e_rsci_idat[234:230]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0
      = conv_s2s_5_6(delay_lane_e_47_sva) + conv_s2s_5_6(taps_e_rsci_idat[239:235]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0
      = conv_s2s_5_6(delay_lane_e_48_sva) + conv_s2s_5_6(taps_e_rsci_idat[244:240]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0
      = conv_s2s_5_6(delay_lane_e_3_sva) + conv_s2s_5_6(taps_e_rsci_idat[19:15]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0
      = conv_s2s_5_6(delay_lane_e_49_sva) + conv_s2s_5_6(taps_e_rsci_idat[249:245]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0
      = conv_s2s_5_6(delay_lane_e_50_sva) + conv_s2s_5_6(taps_e_rsci_idat[254:250]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0
      = conv_s2s_5_6(delay_lane_e_51_sva) + conv_s2s_5_6(taps_e_rsci_idat[259:255]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0
      = conv_s2s_5_6(delay_lane_e_52_sva) + conv_s2s_5_6(taps_e_rsci_idat[264:260]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0
      = conv_s2s_5_6(delay_lane_e_53_sva) + conv_s2s_5_6(taps_e_rsci_idat[269:265]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0
      = conv_s2s_5_6(delay_lane_e_54_sva) + conv_s2s_5_6(taps_e_rsci_idat[274:270]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0
      = conv_s2s_5_6(delay_lane_e_55_sva) + conv_s2s_5_6(taps_e_rsci_idat[279:275]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0
      = conv_s2s_5_6(delay_lane_e_56_sva) + conv_s2s_5_6(taps_e_rsci_idat[284:280]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0
      = conv_s2s_5_6(delay_lane_e_57_sva) + conv_s2s_5_6(taps_e_rsci_idat[289:285]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0
      = conv_s2s_5_6(delay_lane_e_58_sva) + conv_s2s_5_6(taps_e_rsci_idat[294:290]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0
      = conv_s2s_5_6(delay_lane_e_4_sva) + conv_s2s_5_6(taps_e_rsci_idat[24:20]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0
      = conv_s2s_5_6(delay_lane_e_59_sva) + conv_s2s_5_6(taps_e_rsci_idat[299:295]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0
      = conv_s2s_5_6(delay_lane_e_60_sva) + conv_s2s_5_6(taps_e_rsci_idat[304:300]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0
      = conv_s2s_5_6(delay_lane_e_61_sva) + conv_s2s_5_6(taps_e_rsci_idat[309:305]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0
      = conv_s2s_5_6(delay_lane_e_62_sva) + conv_s2s_5_6(taps_e_rsci_idat[314:310]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0
      = conv_s2s_5_6({MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      , MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1})
      + conv_s2s_5_6(taps_e_rsci_idat[319:315]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0
      = conv_s2s_5_6(delay_lane_e_5_sva) + conv_s2s_5_6(taps_e_rsci_idat[29:25]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0
      = conv_s2s_5_6(delay_lane_e_6_sva) + conv_s2s_5_6(taps_e_rsci_idat[34:30]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0
      = conv_s2s_5_6(delay_lane_e_7_sva) + conv_s2s_5_6(taps_e_rsci_idat[39:35]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0[5:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0
      = conv_s2s_5_6(delay_lane_e_8_sva) + conv_s2s_5_6(taps_e_rsci_idat[44:40]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0 =
      nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0[5:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc = and_dcpl_109
      | and_dcpl_154 | and_dcpl_157;
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= 22'b0000000000000000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_e_rsci_idat <= 5'b00000;
    end
    else if ( (and_dcpl_86 & (~ (fsm_output[3])) & and_dcpl_85 & (fsm_output[0])
        & (~ (fsm_output[6])) & (~ (fsm_output[2])) & or_dcpl_105) | return_e_rsci_idat_mx0c1
        ) begin
      return_e_rsci_idat <= MUX_v_5_2_2((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[4:0]),
          5'b01111, return_e_rsci_idat_mx0c1);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      return_m_rsci_idat <= 11'b00000000000;
    end
    else if ( ~((~ (fsm_output[8])) | (fsm_output[1]) | (~ (fsm_output[0])) | or_dcpl_99
        | or_dcpl_98) ) begin
      return_m_rsci_idat <= MUX1HOT_v_11_3_2(11'b01111111111, 11'b10000000000, (MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:2]),
          {result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_63_nl
          , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_or_cse
        ) begin
      MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl,
          and_dcpl_109);
      MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl,
          and_dcpl_109);
      MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl,
          and_dcpl_109);
      MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl,
          and_dcpl_109);
      MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl,
          and_dcpl_109);
      MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl,
          and_dcpl_109);
      MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl,
          and_dcpl_109);
      MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl,
          and_dcpl_109);
      MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl,
          and_dcpl_109);
      MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl,
          and_dcpl_109);
      MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl,
          and_dcpl_109);
      MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl,
          and_dcpl_109);
      MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl,
          and_dcpl_109);
      MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl,
          and_dcpl_109);
      MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= MUX_s_1_2_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_14_nl,
          and_dcpl_109);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= 1'b0;
    end
    else if ( ~ or_dcpl_103 ) begin
      MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm
          <= ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[3:0]!=4'b0000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_64_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_63_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_62_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_61_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_60_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_59_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_58_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_57_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_56_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_55_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_54_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_53_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_52_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_51_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_50_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_49_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_48_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_47_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_46_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_45_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_44_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_43_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_42_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_41_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_40_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_39_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_38_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_37_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_36_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_35_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_34_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_33_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= 1'b0;
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= 1'b0;
      reg_return_e_triosy_obj_ld_cse <= 1'b0;
      reg_taps_e_triosy_obj_ld_cse <= 1'b0;
      MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= 18'b000000000000000000;
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= 18'b000000000000000000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva <=
          4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1
          <= 2'b00;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm
          <= 4'b0000;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1
          <= 2'b00;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0 <=
          1'b0;
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1 <=
          4'b0000;
    end
    else begin
      MAC_64_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0!=22'b0000000000000000000000);
      MAC_63_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0!=22'b0000000000000000000000);
      MAC_62_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0!=22'b0000000000000000000000);
      MAC_61_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0!=22'b0000000000000000000000);
      MAC_60_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0!=22'b0000000000000000000000);
      MAC_59_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0!=22'b0000000000000000000000);
      MAC_58_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0!=22'b0000000000000000000000);
      MAC_57_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0!=22'b0000000000000000000000);
      MAC_56_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0!=22'b0000000000000000000000);
      MAC_55_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0!=22'b0000000000000000000000);
      MAC_54_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0!=22'b0000000000000000000000);
      MAC_53_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0!=22'b0000000000000000000000);
      MAC_52_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0!=22'b0000000000000000000000);
      MAC_51_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0!=22'b0000000000000000000000);
      MAC_50_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0!=22'b0000000000000000000000);
      MAC_49_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0!=22'b0000000000000000000000);
      MAC_48_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0!=22'b0000000000000000000000);
      MAC_47_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0!=22'b0000000000000000000000);
      MAC_46_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0!=22'b0000000000000000000000);
      MAC_45_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0!=22'b0000000000000000000000);
      MAC_44_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0!=22'b0000000000000000000000);
      MAC_43_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0!=22'b0000000000000000000000);
      MAC_42_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0!=22'b0000000000000000000000);
      MAC_41_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0!=22'b0000000000000000000000);
      MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_40_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0!=22'b0000000000000000000000);
      MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_39_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0!=22'b0000000000000000000000);
      MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_38_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0!=22'b0000000000000000000000);
      MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_37_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0!=22'b0000000000000000000000);
      MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_36_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0!=22'b0000000000000000000000);
      MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_35_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0!=22'b0000000000000000000000);
      MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_34_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0!=22'b0000000000000000000000);
      MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_33_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0!=22'b0000000000000000000000);
      MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0!=22'b0000000000000000000000);
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0!=22'b0000000000000000000000);
      MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0!=22'b0000000000000000000000);
      MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0!=22'b0000000000000000000000);
      MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0!=22'b0000000000000000000000);
      MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0!=22'b0000000000000000000000);
      MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0!=22'b0000000000000000000000);
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0!=22'b0000000000000000000000);
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0!=22'b0000000000000000000000);
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_15_nl,
          and_dcpl_109);
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_16_nl,
          and_dcpl_109);
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_17_nl,
          and_dcpl_109);
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_18_nl,
          and_dcpl_109);
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_19_nl,
          and_dcpl_109);
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_20_nl,
          and_dcpl_109);
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_21_nl,
          and_dcpl_109);
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_22_nl,
          and_dcpl_109);
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_23_nl,
          and_dcpl_109);
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_24_nl,
          and_dcpl_109);
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_25_nl,
          and_dcpl_109);
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_26_nl,
          and_dcpl_109);
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_27_nl,
          and_dcpl_109);
      MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_28_nl,
          and_dcpl_109);
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0!=22'b0000000000000000000000);
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0!=22'b0000000000000000000000);
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0!=22'b0000000000000000000000);
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0!=22'b0000000000000000000000);
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0!=22'b0000000000000000000000);
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0!=22'b0000000000000000000000);
      MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0!=22'b0000000000000000000000);
      MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0!=22'b0000000000000000000000);
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5 <= MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[5];
      MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm <= MUX_s_1_2_2(MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_29_nl,
          and_dcpl_109);
      reg_return_e_triosy_obj_ld_cse <= and_dcpl_97 & and_dcpl_95 & and_dcpl_101;
      reg_taps_e_triosy_obj_ld_cse <= ~ or_dcpl_103;
      MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_34_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_35_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_36_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_37_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_38_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_39_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_40_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_41_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_42_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_43_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_44_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_45_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_46_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_47_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_48_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_49_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_50_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_51_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_52_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_53_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_54_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_55_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_56_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_57_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_58_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_59_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_60_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_61_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_62_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_63_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_sva_mx0w0[21:4];
      MAC_1_leading_sign_18_1_1_0_cmp_mantissa <= ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[21:4];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_124_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_120_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_116_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_96_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6
          <= MUX_s_1_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1[6]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
          <= MUX1HOT_s_1_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0[5]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1[5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5
          <= MUX_v_2_2_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:5]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl,
          and_dcpl_109);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_10_itm
          <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg[3:0]),
          (z_out_1[3:0]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]),
          (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
          {and_251_nl , and_254_nl , and_257_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_4_sva_2_1
          <= MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_13_itm
          <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg[3:0]),
          MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_56, leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_57,
          {and_261_nl , and_264_nl , and_267_nl , and_dcpl_151 , and_dcpl_245});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_5_sva_2_1
          <= MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_6_sva_2_1
          <= MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_7_sva_2_1
          <= MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_22_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[3:0]),
          MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_43_nl , and_274_nl , (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_8_sva_2_1
          <= MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_25_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg[3:0]),
          MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_44_nl , and_276_nl , (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_9_sva_2_1
          <= MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_10_sva <=
          MUX1HOT_v_4_4_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[3:0]), (z_out[3:0]), {and_279_nl
          , and_284_nl , and_287_nl , and_dcpl_151});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_10_sva_2_1
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_31_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg[3:0]),
          MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_27_nl , and_289_nl , (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_11_sva_2_1
          <= MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_34_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg[3:0]),
          MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_28_nl , and_291_nl , (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_12_sva_2_1
          <= MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_37_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg[3:0]),
          MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_29_nl , and_293_nl , (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_13_sva_2_1
          <= MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_40_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[3:0]),
          MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_30_nl , and_295_nl , (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_14_sva_2_1
          <= MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_43_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg[3:0]),
          MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_31_nl , and_297_nl , (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_15_sva_2_1
          <= MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_46_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg[3:0]),
          MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_32_nl , and_299_nl , (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_16_sva_2_1
          <= MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_49_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg[3:0]),
          MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_33_nl , and_301_nl , (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_17_sva_2_1
          <= MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_52_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[3:0]),
          MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_34_nl , and_303_nl , (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_18_sva_2_1
          <= MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_55_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg[3:0]),
          MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_35_nl , and_305_nl , (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_19_sva_2_1
          <= MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_58_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg[3:0]),
          MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_36_nl , and_307_nl , (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_20_sva_2_1
          <= MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_61_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[3:0]),
          MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_37_nl , and_309_nl , (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_21_sva_2_1
          <= MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_64_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[3:0]),
          MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_39_nl , and_311_nl , (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_22_sva_2_1
          <= MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_67_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[3:0]),
          MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_40_nl , and_313_nl , (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_23_sva_2_1
          <= MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_70_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[3:0]),
          MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_298_nl , and_315_nl , (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_24_sva_2_1
          <= MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_73_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[3:0]),
          MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_299_nl , and_317_nl , (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_25_sva_2_1
          <= MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_76_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[3:0]),
          MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_300_nl , and_319_nl , (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_26_sva_2_1
          <= MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_79_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[3:0]),
          MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_301_nl , and_321_nl , (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_27_sva_2_1
          <= MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_82_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[3:0]),
          MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_302_nl , and_323_nl , (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_28_sva_2_1
          <= MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_85_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[3:0]),
          MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_303_nl , and_325_nl , (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_29_sva_2_1
          <= MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_88_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[3:0]),
          MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_304_nl , and_327_nl , (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_30_sva_2_1
          <= MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_91_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[3:0]),
          MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_305_nl , and_329_nl , (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_31_sva_2_1
          <= MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_94_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[3:0]),
          MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_306_nl , and_331_nl , (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_32_sva_2_1
          <= MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_97_itm
          <= MUX1HOT_v_4_3_2((MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg[3:0]),
          MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          {nor_307_nl , and_333_nl , (MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])});
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_33_sva_2_1
          <= MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0 <=
          MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl,
          (MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4]), mux_194_itm);
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1 <=
          MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl,
          (MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[3:0]),
          mux_194_itm);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_770_rgt | and_930_rgt ) begin
      MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0,
          {(~ and_118_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl
          , and_930_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_756_rgt | and_922_rgt ) begin
      MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0,
          {(~ and_119_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl
          , and_922_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_749_rgt | and_918_rgt ) begin
      MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0,
          {(~ and_120_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl
          , and_918_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_743_rgt | and_913_rgt ) begin
      MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0,
          {(~ and_121_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl
          , and_913_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_737_rgt | and_909_rgt ) begin
      MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0,
          {(~ and_122_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl
          , and_909_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_729_rgt | and_905_rgt ) begin
      MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_33_lpi_1_dfm_1[4:0]),
          {(~ nor_248_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl
          , and_905_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_723_rgt | and_901_rgt ) begin
      MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_32_lpi_1_dfm_1[4:0]),
          {(~ and_125_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl
          , and_901_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_717_rgt | and_897_rgt ) begin
      MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_31_lpi_1_dfm_1[4:0]),
          {(~ and_127_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl
          , and_897_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_710_rgt | and_893_rgt ) begin
      MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_30_lpi_1_dfm_1[4:0]),
          {(~ and_129_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl
          , and_893_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_704_rgt | and_890_rgt ) begin
      MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_62_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_3_lpi_1_dfm_1[4:0]),
          {(~ and_133_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl
          , and_890_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_697_rgt | and_884_rgt ) begin
      MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_29_lpi_1_dfm_1[4:0]),
          {(~ and_135_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl
          , and_884_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_683_rgt | and_876_rgt ) begin
      MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_27_lpi_1_dfm_1[4:0]),
          {(~ and_137_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl
          , and_876_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_675_rgt | and_872_rgt ) begin
      MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_26_lpi_1_dfm_1[4:0]),
          {(~ and_138_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl
          , and_872_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_667_rgt | and_868_rgt ) begin
      MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_25_lpi_1_dfm_1[4:0]),
          {(~ and_139_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl
          , and_868_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_660_rgt | and_864_rgt ) begin
      MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_24_lpi_1_dfm_1[4:0]),
          {(~ and_140_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl
          , and_864_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_653_rgt | and_860_rgt ) begin
      MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_23_lpi_1_dfm_1[4:0]),
          {(~ and_141_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_46_nl
          , and_860_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_646_rgt | and_856_rgt ) begin
      MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_22_lpi_1_dfm_1[4:0]),
          {(~ and_142_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_49_nl
          , and_856_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_639_rgt | and_852_rgt ) begin
      MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_21_lpi_1_dfm_1[4:0]),
          {(~ and_143_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_52_nl
          , and_852_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_631_rgt | and_848_rgt ) begin
      MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_20_lpi_1_dfm_1[4:0]),
          {(~ and_144_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_55_nl
          , and_848_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_470_rgt | and_559_rgt ) begin
      MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_19_lpi_1_dfm_1[4:0]),
          {(~ and_145_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_58_nl
          , and_559_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_453_rgt | and_551_rgt ) begin
      MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_17_lpi_1_dfm_1[4:0]),
          {(~ and_146_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_61_nl
          , and_551_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_445_rgt | and_547_rgt ) begin
      MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_16_lpi_1_dfm_1[4:0]),
          {(~ and_149_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_64_nl
          , and_547_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_437_rgt | and_543_rgt ) begin
      MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_15_lpi_1_dfm_1[4:0]),
          {(~ and_151_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_67_nl
          , and_543_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_430_rgt | and_539_rgt ) begin
      MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_14_lpi_1_dfm_1[4:0]),
          {(~ and_153_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_70_nl
          , and_539_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_422_rgt | and_535_rgt ) begin
      MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_13_lpi_1_dfm_1[4:0]),
          {(~ and_155_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_73_nl
          , and_535_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_415_rgt | and_531_rgt ) begin
      MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_12_lpi_1_dfm_1[4:0]),
          {(~ and_156_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_76_nl
          , and_531_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_408_rgt | and_527_rgt ) begin
      MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_11_lpi_1_dfm_1[4:0]),
          {(~ and_158_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_79_nl
          , and_527_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_401_rgt | and_523_rgt ) begin
      MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_10_lpi_1_dfm_1[4:0]),
          {(~ and_159_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_82_nl
          , and_523_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_763_rgt | and_926_rgt ) begin
      MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg, 5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0,
          {(~ and_160_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_85_nl
          , and_926_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_690_rgt | and_880_rgt ) begin
      MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_28_lpi_1_dfm_1[4:0]),
          {(~ and_161_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_88_nl
          , and_880_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= 5'b00000;
    end
    else if ( and_dcpl_109 | or_462_rgt | and_555_rgt ) begin
      MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0 <= MUX1HOT_v_5_4_2((MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm[4:0]),
          MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg, 5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_18_lpi_1_dfm_1[4:0]),
          {(~ and_162_rgt) , and_dcpl_109 , ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_91_nl
          , and_555_rgt});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_1_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_103 ) begin
      delay_lane_e_1_sva <= delay_lane_e_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_1_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      delay_lane_m_1_sva <= delay_lane_m_0_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_0_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_103 ) begin
      delay_lane_e_0_sva <= input_e_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_0_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_103 ) begin
      delay_lane_m_0_sva <= input_m_rsci_idat;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_62_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_62_sva <= delay_lane_e_61_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_62_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_62_sva <= delay_lane_m_61_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_61_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_61_sva <= delay_lane_e_60_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_61_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_61_sva <= delay_lane_m_60_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_60_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_60_sva <= delay_lane_e_59_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_60_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_60_sva <= delay_lane_m_59_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_59_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_59_sva <= delay_lane_e_58_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_59_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_59_sva <= delay_lane_m_58_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_58_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_58_sva <= delay_lane_e_57_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_58_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_58_sva <= delay_lane_m_57_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_57_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_57_sva <= delay_lane_e_56_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_57_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_57_sva <= delay_lane_m_56_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_56_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_56_sva <= delay_lane_e_55_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_56_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_56_sva <= delay_lane_m_55_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_55_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_55_sva <= delay_lane_e_54_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_55_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_55_sva <= delay_lane_m_54_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_54_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_54_sva <= delay_lane_e_53_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_54_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_54_sva <= delay_lane_m_53_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_53_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_53_sva <= delay_lane_e_52_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_53_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_53_sva <= delay_lane_m_52_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_52_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_52_sva <= delay_lane_e_51_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_52_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_52_sva <= delay_lane_m_51_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_51_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_51_sva <= delay_lane_e_50_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_51_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_51_sva <= delay_lane_m_50_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_50_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_50_sva <= delay_lane_e_49_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_50_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_50_sva <= delay_lane_m_49_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_49_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_49_sva <= delay_lane_e_48_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_49_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_49_sva <= delay_lane_m_48_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_48_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_48_sva <= delay_lane_e_47_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_48_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_48_sva <= delay_lane_m_47_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_47_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_47_sva <= delay_lane_e_46_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_47_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_47_sva <= delay_lane_m_46_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_46_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_46_sva <= delay_lane_e_45_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_46_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_46_sva <= delay_lane_m_45_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_45_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_45_sva <= delay_lane_e_44_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_45_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_45_sva <= delay_lane_m_44_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_44_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_44_sva <= delay_lane_e_43_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_44_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_44_sva <= delay_lane_m_43_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_43_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_43_sva <= delay_lane_e_42_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_43_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_43_sva <= delay_lane_m_42_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_42_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_42_sva <= delay_lane_e_41_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_42_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_42_sva <= delay_lane_m_41_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_41_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_41_sva <= delay_lane_e_40_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_41_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_41_sva <= delay_lane_m_40_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_40_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_40_sva <= delay_lane_e_39_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_40_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_40_sva <= delay_lane_m_39_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_39_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_39_sva <= delay_lane_e_38_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_39_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_39_sva <= delay_lane_m_38_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_38_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_38_sva <= delay_lane_e_37_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_38_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_38_sva <= delay_lane_m_37_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_37_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_37_sva <= delay_lane_e_36_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_37_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_37_sva <= delay_lane_m_36_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_36_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_36_sva <= delay_lane_e_35_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_36_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_36_sva <= delay_lane_m_35_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_35_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_35_sva <= delay_lane_e_34_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_35_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_35_sva <= delay_lane_m_34_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_34_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_34_sva <= delay_lane_e_33_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_34_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_34_sva <= delay_lane_m_33_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_33_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_33_sva <= delay_lane_e_32_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_33_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_33_sva <= delay_lane_m_32_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_32_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_32_sva <= delay_lane_e_31_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_32_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_32_sva <= delay_lane_m_31_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_31_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_31_sva <= delay_lane_e_30_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_31_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_31_sva <= delay_lane_m_30_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_30_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_30_sva <= delay_lane_e_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_30_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_30_sva <= delay_lane_m_29_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_29_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_29_sva <= delay_lane_e_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_29_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_29_sva <= delay_lane_m_28_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_28_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_28_sva <= delay_lane_e_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_28_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_28_sva <= delay_lane_m_27_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_27_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_27_sva <= delay_lane_e_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_27_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_27_sva <= delay_lane_m_26_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_26_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_26_sva <= delay_lane_e_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_26_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_26_sva <= delay_lane_m_25_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_25_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_25_sva <= delay_lane_e_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_25_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_25_sva <= delay_lane_m_24_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_24_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_24_sva <= delay_lane_e_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_24_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_24_sva <= delay_lane_m_23_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_23_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_23_sva <= delay_lane_e_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_23_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_23_sva <= delay_lane_m_22_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_22_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_22_sva <= delay_lane_e_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_22_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_22_sva <= delay_lane_m_21_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_21_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_21_sva <= delay_lane_e_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_21_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_21_sva <= delay_lane_m_20_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_20_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_20_sva <= delay_lane_e_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_20_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_20_sva <= delay_lane_m_19_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_19_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_19_sva <= delay_lane_e_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_19_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_19_sva <= delay_lane_m_18_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_18_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_18_sva <= delay_lane_e_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_18_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_18_sva <= delay_lane_m_17_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_17_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_17_sva <= delay_lane_e_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_17_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_17_sva <= delay_lane_m_16_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_16_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_16_sva <= delay_lane_e_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_16_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_16_sva <= delay_lane_m_15_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_15_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_15_sva <= delay_lane_e_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_15_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_15_sva <= delay_lane_m_14_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_14_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_14_sva <= delay_lane_e_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_14_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_14_sva <= delay_lane_m_13_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_13_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_13_sva <= delay_lane_e_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_13_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_13_sva <= delay_lane_m_12_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_12_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_12_sva <= delay_lane_e_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_12_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_12_sva <= delay_lane_m_11_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_11_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_11_sva <= delay_lane_e_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_11_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_11_sva <= delay_lane_m_10_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_10_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_10_sva <= delay_lane_e_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_10_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_10_sva <= delay_lane_m_9_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_9_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_9_sva <= delay_lane_e_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_9_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_9_sva <= delay_lane_m_8_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_8_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_8_sva <= delay_lane_e_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_8_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_8_sva <= delay_lane_m_7_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_7_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_7_sva <= delay_lane_e_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_7_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_7_sva <= delay_lane_m_6_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_6_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_6_sva <= delay_lane_e_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_6_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_6_sva <= delay_lane_m_5_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_5_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_5_sva <= delay_lane_e_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_5_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_5_sva <= delay_lane_m_4_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_4_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_4_sva <= delay_lane_e_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_4_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_4_sva <= delay_lane_m_3_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_3_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_3_sva <= delay_lane_e_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_3_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_3_sva <= delay_lane_m_2_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_e_2_sva <= 5'b00000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_e_2_sva <= delay_lane_e_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      delay_lane_m_2_sva <= 11'b00000000000;
    end
    else if ( ~ or_dcpl_120 ) begin
      delay_lane_m_2_sva <= delay_lane_m_1_sva;
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
          <= 1'b0;
    end
    else if ( and_dcpl_105 | and_dcpl_109 | and_dcpl_151 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm
          <= MUX1HOT_s_1_5_2(MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl,
          (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_60_rtn_oreg[4]), (MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
          (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
          {and_dcpl_105 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_2_cse
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_3_cse});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7 <= 4'b0000;
    end
    else if ( ~(mux_1109_nl | (fsm_output[8])) ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_10_7 <= MUX1HOT_v_4_128_2((MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]),
          result_m_1_lpi_1_dfm_1_10_7, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_10_7,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10:7]),
          (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10:7]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7,
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7,
          (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7,
          (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7,
          (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7,
          (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[10:7]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[10:7]),
          (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[10:7]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[10:7]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[10:7]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[10:7]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[10:7]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[10:7]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[10:7]),
          (MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[10:7]),
          (MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[10:7]),
          (MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[10:7]),
          (MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[10:7]),
          (MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[10:7]),
          (MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[10:7]),
          (MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[10:7]),
          (MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[10:7]),
          (MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[10:7]),
          (MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[10:7]),
          (MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[10:7]),
          (MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[10:7]),
          (MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[10:7]),
          (MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[10:7]),
          (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[10:7]),
          (MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[10:7]),
          (MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[10:7]),
          (MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[10:7]),
          (MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[10:7]),
          (MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[10:7]),
          (MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[10:7]),
          (MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7,
          (MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_41_lpi_1_dfm_10_7,
          (MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_42_lpi_1_dfm_10_7,
          (MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_43_lpi_1_dfm_10_7,
          (MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_44_lpi_1_dfm_10_7,
          (MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_45_lpi_1_dfm_10_7,
          (MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_46_lpi_1_dfm_10_7,
          (MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_47_lpi_1_dfm_10_7,
          (MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_48_lpi_1_dfm_10_7,
          (MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_49_lpi_1_dfm_10_7,
          (MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_50_lpi_1_dfm_10_7,
          (MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_51_lpi_1_dfm_10_7,
          (MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_52_lpi_1_dfm_10_7,
          (MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_53_lpi_1_dfm_10_7,
          (MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_54_lpi_1_dfm_10_7,
          (MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_55_lpi_1_dfm_10_7,
          (MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_56_lpi_1_dfm_10_7,
          (MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_57_lpi_1_dfm_10_7,
          (MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_58_lpi_1_dfm_10_7,
          (MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_59_lpi_1_dfm_10_7,
          (MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_60_lpi_1_dfm_10_7,
          (MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_61_lpi_1_dfm_10_7,
          (MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_62_lpi_1_dfm_10_7,
          (MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_63_lpi_1_dfm_10_7,
          (MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12:9]), MAC_ac_float_cctor_m_lpi_1_dfm_10_7,
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[10:7]), {and_dcpl_221
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse
          , and_dcpl_157});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(mux_657_nl & and_184_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_417_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_4_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_312_nl
          , and_1301_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_639_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_419_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_310_nl
          , and_1277_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_635_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_421_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_92_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_308_nl
          , and_1273_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_632_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_423_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_306_nl
          , and_1269_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_629_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_425_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_304_nl
          , and_1265_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_626_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_427_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_302_nl
          , and_1261_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_621_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_429_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_300_nl
          , and_1257_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_618_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_431_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_298_nl
          , and_1253_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_615_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_433_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_296_nl
          , and_1249_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_611_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_435_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_294_nl
          , and_1244_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_608_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_437_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_292_nl
          , and_1240_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_654_nl) & and_196_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_439_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_5_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_291_nl
          , and_1297_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_604_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_441_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_289_nl
          , and_1235_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_601_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_443_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_287_nl
          , and_1231_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_598_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_445_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_285_nl
          , and_1227_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_594_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_447_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_283_nl
          , and_1223_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_591_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_449_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_281_nl
          , and_1219_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_588_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_451_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_279_nl
          , and_1215_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_584_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_453_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_277_nl
          , and_1210_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_582_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_455_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_275_nl
          , and_1206_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_578_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_457_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_273_nl
          , and_1201_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_576_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_459_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_271_nl
          , and_1197_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_651_nl) & and_210_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_461_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_6_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_270_nl
          , and_1293_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_574_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_463_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_268_nl
          , and_1193_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_570_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_465_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_266_nl
          , and_1189_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_568_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_467_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_264_nl
          , and_1185_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( mux_566_nl | (fsm_output[8]) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_469_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl,
          5'b01111, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0,
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_262_nl
          , and_1181_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_648_nl) & and_219_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_471_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_7_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_261_nl
          , and_1289_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_645_nl) & and_220_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_473_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_8_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_260_nl
          , and_1285_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~((~ mux_642_nl) & and_221_ssc) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_5_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_conc_475_itm_5_0[4:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl,
          5'b01111, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_9_lpi_1_dfm_1[4:0]),
          {and_dcpl_105 , and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_259_nl
          , and_1281_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 3'b000;
    end
    else if ( and_dcpl_160 | and_dcpl_151 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= MUX_v_3_2_2(MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp,
          and_dcpl_151);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= 3'b000;
    end
    else if ( ~ or_dcpl_134 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
          <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva <= 7'b0000000;
    end
    else if ( ~(mux_260_nl & and_dcpl_1 & and_dcpl_101) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva <= nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[6:0];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= 5'b00000;
    end
    else if ( ~(((nor_518_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_6_5[1]))
        & and_dcpl_152 & and_dcpl_497) | (~(mux_559_nl | (fsm_output[8])))) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0
          <= MUX1HOT_v_5_3_2((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[4:0]),
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_64_nl,
          5'b01111, {and_dcpl_160 , and_dcpl_109 , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc ) begin
      MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7 <= MUX_v_4_2_2((z_out_2[10:7]), (delay_lane_m_62_sva[10:7]),
          and_dcpl_207);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_ssc & (~ and_dcpl_109) ) begin
      MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0 <= MUX1HOT_v_7_3_2(MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (z_out_2[6:0]), (delay_lane_m_62_sva[6:0]), {and_dcpl_203 , and_dcpl_154
          , and_dcpl_207});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_41_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_42_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_43_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_44_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_45_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_46_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_47_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_48_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_49_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_50_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_51_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_52_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_53_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_54_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_55_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_56_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_57_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_58_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_59_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_60_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_61_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_62_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_63_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7 <= 4'b0000;
      MAC_ac_float_cctor_m_lpi_1_dfm_10_7 <= 4'b0000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_or_1_cse ) begin
      MAC_ac_float_cctor_m_41_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_41_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_42_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_42_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_43_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_43_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_44_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_44_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_45_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_45_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_46_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_46_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_47_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_47_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_48_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_48_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_49_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_49_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_50_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_50_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_51_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_51_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_52_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_52_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_53_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_53_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_54_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_54_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_55_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_55_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_56_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_56_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_57_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_57_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_58_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_58_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_59_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_59_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_60_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_60_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_61_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_61_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_62_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_62_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_63_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_63_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1[10:7];
      MAC_ac_float_cctor_m_lpi_1_dfm_10_7 <= MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1[10:7];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 <= 7'b0000000;
      MAC_ac_float_cctor_m_lpi_1_dfm_6_0 <= 7'b0000000;
    end
    else if ( ac_float_cctor_ac_float_22_2_6_AC_TRN_and_1_cse ) begin
      MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_41_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_42_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_43_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_44_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_45_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_46_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_47_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_48_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_49_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_50_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_51_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_52_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_53_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_54_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_55_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_56_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_57_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_58_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_59_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_60_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_61_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_62_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_63_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
      MAC_ac_float_cctor_m_lpi_1_dfm_6_0 <= MUX_v_7_2_2(MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl,
          (MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1[6:0]), and_dcpl_154);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
        | and_dcpl_221 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva <= MUX1HOT_v_11_5_2((MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_1_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), (MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_2_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c1
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c2
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva_mx0c3
          , and_dcpl_221});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
          <= 1'b0;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_or_cse
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_2_sva
          <= MUX_s_1_2_2((~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_4_sva
          <= MUX_s_1_2_2((~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_33_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_5_sva
          <= MUX_s_1_2_2((~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_34_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_6_sva
          <= MUX_s_1_2_2((~ MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_35_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_7_sva
          <= MUX_s_1_2_2((~ MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_36_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_8_sva
          <= MUX_s_1_2_2((~ MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_37_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_9_sva
          <= MUX_s_1_2_2((~ MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_38_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_12_sva
          <= MUX_s_1_2_2((~ MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_13_sva
          <= MUX_s_1_2_2((~ MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_14_sva
          <= MUX_s_1_2_2((~ MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_15_sva
          <= MUX_s_1_2_2((~ MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_16_sva
          <= MUX_s_1_2_2((~ MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_17_sva
          <= MUX_s_1_2_2((~ MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_18_sva
          <= MUX_s_1_2_2((~ MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_19_sva
          <= MUX_s_1_2_2((~ MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_20_sva
          <= MUX_s_1_2_2((~ MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_21_sva
          <= MUX_s_1_2_2((~ MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_22_sva
          <= MUX_s_1_2_2((~ MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_23_sva
          <= MUX_s_1_2_2((~ MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_24_sva
          <= MUX_s_1_2_2((~ MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_25_sva
          <= MUX_s_1_2_2((~ MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_25_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_26_sva
          <= MUX_s_1_2_2((~ MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_27_sva
          <= MUX_s_1_2_2((~ MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_28_sva
          <= MUX_s_1_2_2((~ MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_29_sva
          <= MUX_s_1_2_2((~ MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_30_sva
          <= MUX_s_1_2_2((~ MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_31_sva
          <= MUX_s_1_2_2((~ MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_32_sva
          <= MUX_s_1_2_2((~ MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_33_sva
          <= MUX_s_1_2_2((~ MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_32_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_nl,
          MAC_59_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_nl,
          MAC_58_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_nl,
          MAC_57_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_nl,
          MAC_55_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_nl,
          MAC_54_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_nl,
          MAC_53_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_nl,
          MAC_52_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_nl,
          MAC_51_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_nl,
          MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_nl,
          MAC_50_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_nl,
          MAC_49_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_nl,
          MAC_48_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_nl,
          MAC_47_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_nl,
          MAC_46_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_nl,
          MAC_45_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_nl,
          MAC_44_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl,
          MAC_43_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl,
          MAC_42_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl,
          MAC_41_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl,
          MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl,
          MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl,
          MAC_39_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl,
          ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_nl,
          and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl,
          MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl,
          MAC_63_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl,
          MAC_62_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl,
          MAC_61_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl,
          MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl,
          MAC_60_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
          <= MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl,
          MAC_56_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, and_dcpl_154);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
          <= MUX_s_1_2_2(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same_oreg, MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl,
          and_dcpl_154);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1
          <= 2'b00;
    end
    else if ( ~(or_151_cse | or_dcpl_99 | or_dcpl_98) ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_2_sva_2_1
          <= MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2:1];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= 1'b0;
    end
    else if ( and_dcpl_109 | and_dcpl_151 | and_dcpl_221 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_10_sva
          <= MUX1HOT_s_1_3_2((~ MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          (~ MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl, {and_dcpl_109
          , and_dcpl_151 , and_dcpl_221});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= 1'b0;
    end
    else if ( and_dcpl_109 | and_dcpl_151 | and_dcpl_245 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva
          <= MUX1HOT_s_1_3_2((~ MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1),
          MAC_2_ac_float_cctor_operator_ac_float_cctor_operator_nor_cse, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_51_nl,
          {and_dcpl_109 , and_dcpl_151 , and_dcpl_245});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva <= MUX1HOT_v_11_3_2((MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_34_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva <= MUX1HOT_v_11_3_2((MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_35_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva <= MUX1HOT_v_11_3_2((MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_36_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva <= MUX1HOT_v_11_3_2((MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_37_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva <= MUX1HOT_v_11_3_2((MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_38_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva <= MUX1HOT_v_11_3_2((MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_39_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva <= MUX1HOT_v_11_3_2((MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_40_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva <= MUX1HOT_v_11_3_2((MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_41_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva <= MUX1HOT_v_11_3_2((MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_42_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva <= MUX1HOT_v_11_3_2((MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_43_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva <= MUX1HOT_v_11_3_2((MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_44_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva <= MUX1HOT_v_11_3_2((MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_45_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva <= MUX1HOT_v_11_3_2((MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_46_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva <= MUX1HOT_v_11_3_2((MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_47_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva <= MUX1HOT_v_11_3_2((MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_48_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva <= MUX1HOT_v_11_3_2((MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_49_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_25_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva <= MUX1HOT_v_11_3_2((MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_50_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva <= MUX1HOT_v_11_3_2((MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_51_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva <= MUX1HOT_v_11_3_2((MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_52_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva <= MUX1HOT_v_11_3_2((MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_53_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva <= MUX1HOT_v_11_3_2((MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_54_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva <= MUX1HOT_v_11_3_2((MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_55_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva <= MUX1HOT_v_11_3_2((MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_56_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_32_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva <= MUX1HOT_v_11_3_2((MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_57_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_33_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva <= MUX1HOT_v_11_3_2((MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_58_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_34_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva <= MUX1HOT_v_11_3_2((MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_59_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_35_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva <= MUX1HOT_v_11_3_2((MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_60_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_36_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva <= MUX1HOT_v_11_3_2((MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_61_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_37_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva <= MUX1HOT_v_11_3_2((MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_62_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_38_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva <= MUX1HOT_v_11_3_2((MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_63_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_39_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva <= 11'b00000000000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
        | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
        | and_dcpl_154 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva <= MUX1HOT_v_11_3_2((MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_rshift_itm[21:11]),
          (MAC_64_operator_22_2_true_AC_TRN_AC_WRAP_lshift_itm[21:11]), MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w2,
          {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c0
          , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva_mx0c1
          , and_dcpl_154});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp <= 1'b0;
    end
    else if ( and_dcpl_109 | and_dcpl_151 | and_dcpl_221 | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3
        ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp <= MUX1HOT_s_1_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl,
          leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_54, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl,
          result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3, {and_dcpl_109
          , and_dcpl_151 , and_dcpl_221 , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_mx0c3});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_10_7 <=
          4'b0000;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_6 <= 1'b0;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_5_4 <=
          2'b00;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0 <=
          4'b0000;
    end
    else if ( result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_ssc ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_10_7 <=
          MUX1HOT_v_4_64_2((z_out_2[10:7]), result_m_1_lpi_1_dfm_1_10_7, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[10:7]),
          MAC_ac_float_cctor_m_5_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_6_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_7_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_8_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_9_lpi_1_dfm_10_7, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[10:7]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[10:7]),
          MAC_ac_float_cctor_m_40_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_41_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_42_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_43_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_44_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_45_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_46_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_47_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_48_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_49_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_50_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_51_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_52_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_53_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_54_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_55_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_56_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_57_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_58_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_59_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_60_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_61_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_62_lpi_1_dfm_10_7, MAC_ac_float_cctor_m_63_lpi_1_dfm_10_7,
          MAC_ac_float_cctor_m_lpi_1_dfm_10_7, {and_dcpl_151 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_6 <= MUX1HOT_s_1_64_2((z_out_2[6]),
          result_m_1_lpi_1_dfm_1_6, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[6]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[6]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[6]),
          (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[6]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[6]),
          (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6]), {and_dcpl_151 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_5_4 <=
          MUX1HOT_v_2_64_2((z_out_2[5:4]), result_m_1_lpi_1_dfm_1_5_4, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[5:4]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[5:4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[5:4]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[5:4]),
          (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[5:4]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[5:4]),
          (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[5:4]), {and_dcpl_151 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64});
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0 <=
          MUX1HOT_v_4_66_2((MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]), (MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg[3:0]),
          MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (z_out_2[3:0]), result_m_1_lpi_1_dfm_1_3_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[3:0]),
          (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[3:0]),
          (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[3:0]),
          (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[3:0]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[3:0]),
          (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]), {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl
          , and_270_nl , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl
          , and_dcpl_151 , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c2
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c3
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c4
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c5
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c6
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c8
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c9
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c10
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c11
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c12
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c13
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c14
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c15
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c16
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c17
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c18
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c19
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c20
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c21
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c22
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c23
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c24
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c25
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c26
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c27
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c28
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c29
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c30
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c31
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c32
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c33
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c34
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c35
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c36
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c37
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c38
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c39
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c40
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c41
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c42
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c43
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c44
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c45
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c46
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c47
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c48
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c49
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c50
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c51
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c52
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c53
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c54
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c55
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c56
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c57
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c58
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c59
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c60
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c61
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c62
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c63
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c64});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_316 ) begin
      ac_float_cctor_operator_return_sva <= ~((MAC_ac_float_cctor_m_lpi_1_dfm_mx0w1!=11'b00000000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_operator_return_9_sva <= 1'b0;
    end
    else if ( ~ or_dcpl_316 ) begin
      ac_float_cctor_operator_return_9_sva <= ~((MAC_ac_float_cctor_m_10_lpi_1_dfm_mx0w2!=11'b00000000000));
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= 2'b00;
    end
    else if ( and_dcpl_154 | and_dcpl_157 ) begin
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_1_sva
          <= MUX_v_2_2_2(MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl,
          and_dcpl_157);
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
          <= 1'b0;
    end
    else if ( ~ and_dcpl_109 ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_0
          <= MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[6];
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
          <= 1'b0;
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2
          <= 5'b00000;
    end
    else if ( ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_95_itm
        ) begin
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_1
          <= MUX_s_1_2_2(ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_64_nl,
          (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[5]),
          and_dcpl_160);
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2
          <= MUX1HOT_v_5_5_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[4:0]),
          (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[4:0]),
          (z_out_1[4:0]), (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_itm[4:0]),
          and_1758_nl, {and_dcpl_105 , and_dcpl_154 , and_dcpl_157 , and_dcpl_160
          , and_dcpl_162});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 <= 1'b0;
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1 <= 2'b00;
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 <= 4'b0000;
    end
    else if ( operator_13_2_true_AC_TRN_AC_WRAP_or_ssc ) begin
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_0 <= MUX1HOT_s_1_129_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[6]),
          (MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), result_m_1_lpi_1_dfm_1_6,
          result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_6,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[6]),
          (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[6]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[6]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[6]),
          (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[6]),
          (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[6]),
          (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[6]),
          (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[6]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[6]),
          (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[6]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[6]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[6]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[6]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[6]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[6]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[6]),
          (MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[6]),
          (MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[6]),
          (MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[6]),
          (MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[6]),
          (MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[6]),
          (MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[6]),
          (MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[6]),
          (MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[6]),
          (MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[6]),
          (MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[6]),
          (MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[6]),
          (MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[6]),
          (MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[6]),
          (MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[6]),
          (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[6]),
          (MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[6]),
          (MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[6]),
          (MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[6]),
          (MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[6]),
          (MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[6]),
          (MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[6]),
          (MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[6]),
          (MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[6]),
          (MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[6]),
          (MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[6]),
          (MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[6]),
          (MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[6]),
          (MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[6]),
          (MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[6]),
          (MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[6]),
          (MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[6]),
          (MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[6]),
          (MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[6]),
          (MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[6]),
          (MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[6]),
          (MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[6]),
          (MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[6]),
          (MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[6]),
          (MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[6]),
          (MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[6]),
          (MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[6]),
          (MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[6]),
          (MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[6]),
          (MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[6]),
          (MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[6]),
          (MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[8]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[6]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[6]), {operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1
          , and_dcpl_221 , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse
          , and_dcpl_157});
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1 <= MUX1HOT_v_2_130_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[5:4]),
          (operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[5:4]), (MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]),
          result_m_1_lpi_1_dfm_1_5_4, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_5_4,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[5:4]),
          (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[5:4]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[5:4]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[5:4]),
          (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[5:4]),
          (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[5:4]),
          (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[5:4]),
          (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[5:4]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[5:4]),
          (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[5:4]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[5:4]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[5:4]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[5:4]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[5:4]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[5:4]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[5:4]),
          (MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[5:4]),
          (MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[5:4]),
          (MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[5:4]),
          (MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[5:4]),
          (MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[5:4]),
          (MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[5:4]),
          (MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[5:4]),
          (MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[5:4]),
          (MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[5:4]),
          (MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[5:4]),
          (MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[5:4]),
          (MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[5:4]),
          (MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[5:4]),
          (MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[5:4]),
          (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[5:4]),
          (MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[5:4]),
          (MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[5:4]),
          (MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[5:4]),
          (MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[5:4]),
          (MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[5:4]),
          (MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[5:4]),
          (MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[5:4]),
          (MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[5:4]),
          (MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[5:4]),
          (MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[5:4]),
          (MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[5:4]),
          (MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[5:4]),
          (MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[5:4]),
          (MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[5:4]),
          (MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[5:4]),
          (MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[5:4]),
          (MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[5:4]),
          (MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[5:4]),
          (MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[5:4]),
          (MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[5:4]),
          (MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[5:4]),
          (MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[5:4]),
          (MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[5:4]),
          (MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[5:4]),
          (MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[5:4]),
          (MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[5:4]),
          (MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[5:4]),
          (MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[5:4]),
          (MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[5:4]),
          (MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[5:4]),
          (MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[7:6]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[5:4]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[5:4]), {and_dcpl_105
          , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 , and_dcpl_221
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse
          , and_dcpl_157});
      operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2 <= MUX1HOT_v_4_130_2((operator_13_2_true_AC_TRN_AC_WRAP_conc_2_itm_5_0[3:0]),
          (operator_13_2_true_AC_TRN_AC_WRAP_conc_4_itm_6_0[3:0]), (MAC_1_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]),
          result_m_1_lpi_1_dfm_1_3_0, result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_3_0,
          (MAC_2_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[3:0]),
          (MAC_3_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_sva[3:0]),
          (MAC_4_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]),
          (MAC_5_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]),
          (MAC_6_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]),
          (MAC_7_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]),
          (MAC_8_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]),
          (MAC_9_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_34_sva[3:0]),
          (MAC_10_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_35_sva[3:0]),
          (MAC_11_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_36_sva[3:0]),
          (MAC_12_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_37_sva[3:0]),
          (MAC_13_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_38_sva[3:0]),
          (MAC_14_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_39_sva[3:0]),
          (MAC_15_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[3:0]),
          (MAC_16_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_41_sva[3:0]),
          (MAC_17_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_42_sva[3:0]),
          (MAC_18_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_43_sva[3:0]),
          (MAC_19_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_44_sva[3:0]),
          (MAC_20_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_45_sva[3:0]),
          (MAC_21_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_46_sva[3:0]),
          (MAC_22_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_47_sva[3:0]),
          (MAC_23_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_48_sva[3:0]),
          (MAC_24_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_49_sva[3:0]),
          (MAC_25_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_50_sva[3:0]),
          (MAC_26_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_51_sva[3:0]),
          (MAC_27_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_52_sva[3:0]),
          (MAC_28_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_53_sva[3:0]),
          (MAC_29_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_54_sva[3:0]),
          (MAC_30_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_55_sva[3:0]),
          (MAC_31_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_56_sva[3:0]),
          (MAC_32_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_57_sva[3:0]),
          (MAC_33_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_58_sva[3:0]),
          (MAC_34_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_59_sva[3:0]),
          (MAC_35_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_60_sva[3:0]),
          (MAC_36_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_61_sva[3:0]),
          (MAC_37_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_62_sva[3:0]),
          (MAC_38_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_63_sva[3:0]),
          (MAC_39_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[3:0]),
          (MAC_40_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[3:0]),
          (MAC_41_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[3:0]),
          (MAC_42_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[3:0]),
          (MAC_43_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[3:0]),
          (MAC_44_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[3:0]),
          (MAC_45_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[3:0]),
          (MAC_46_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[3:0]),
          (MAC_47_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[3:0]),
          (MAC_48_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0[3:0]),
          (MAC_49_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[3:0]),
          (MAC_50_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[3:0]),
          (MAC_51_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[3:0]),
          (MAC_52_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[3:0]),
          (MAC_53_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[3:0]),
          (MAC_54_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[3:0]),
          (MAC_55_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[3:0]),
          (MAC_56_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[3:0]),
          (MAC_57_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[3:0]),
          (MAC_58_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[3:0]),
          (MAC_59_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[3:0]),
          (MAC_60_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[3:0]),
          (MAC_61_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[3:0]),
          (MAC_62_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[3:0]),
          (MAC_63_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[5:2]), (MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]),
          (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_6_sva_mx0w3[3:0]), {and_dcpl_105
          , operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_mx0c1 , and_dcpl_221
          , operator_13_2_true_AC_TRN_AC_WRAP_and_1_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_2_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_3_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_4_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_5_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_6_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_7_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_8_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_9_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_10_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_11_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_12_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_13_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_14_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_15_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_16_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_17_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_18_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_19_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_20_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_21_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_22_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_23_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_24_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_25_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_26_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_27_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_28_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_29_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_30_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_31_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_32_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_33_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_34_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_35_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_36_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_37_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_38_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_39_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_40_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_41_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_42_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_43_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_44_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_45_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_46_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_47_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_48_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_49_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_50_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_51_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_52_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_53_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_54_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_55_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_56_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_57_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_58_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_59_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_60_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_61_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_62_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_63_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_64_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_65_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_66_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_67_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_68_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_69_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_70_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_71_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_72_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_73_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_74_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_75_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_76_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_77_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_78_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_79_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_80_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_81_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_82_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_83_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_84_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_85_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_86_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_87_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_88_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_89_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_90_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_91_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_92_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_93_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_94_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_95_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_96_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_97_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_98_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_99_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_100_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_101_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_102_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_103_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_104_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_105_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_106_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_107_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_108_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_109_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_110_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_111_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_112_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_113_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_114_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_115_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_116_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_117_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_118_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_119_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_120_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_121_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_122_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_123_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_124_cse
          , operator_13_2_true_AC_TRN_AC_WRAP_and_125_cse , operator_13_2_true_AC_TRN_AC_WRAP_and_126_cse
          , and_dcpl_157});
    end
  end
  always @(posedge clk) begin
    if ( rst ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0 <= 8'b00000000;
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 <= 4'b0000;
    end
    else if ( result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_or_ssc ) begin
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_0 <= MUX_v_8_2_2((MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:4]),
          (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[11:4]),
          and_dcpl_157);
      result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_12_1_1_sva_rsp_1 <= MUX1HOT_v_4_5_2((MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]),
          (MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg[3:0]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl,
          (MAC_1_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_acc_itm[3:0]),
          {result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl , and_272_nl
          , result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl , and_dcpl_154
          , and_dcpl_157});
    end
  end
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nor_63_nl
      = ~((MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12]) | result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_127_nl = (MAC_64_operator_13_2_true_AC_TRN_AC_WRAP_lshift_itm[12])
      & (~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp_2_mx0w3);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_nl
      = MUX_s_1_2_2((MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_32_rtn_oreg[4]), MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_1_nl
      = MUX_s_1_2_2((MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_34_rtn_oreg[4]), MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_2_nl
      = MUX_s_1_2_2((MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_35_rtn_oreg[4]), MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_3_nl
      = MUX_s_1_2_2((MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_37_rtn_oreg[4]), MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_4_nl
      = MUX_s_1_2_2((MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_39_rtn_oreg[4]), MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_5_nl
      = MUX_s_1_2_2((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_43_rtn_oreg[4]), MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_6_nl
      = MUX_s_1_2_2((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_45_rtn_oreg[4]), MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_7_nl
      = MUX_s_1_2_2((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_47_rtn_oreg[4]), MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_8_nl
      = MUX_s_1_2_2((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_49_rtn_oreg[4]), MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_9_nl
      = MUX_s_1_2_2((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_51_rtn_oreg[4]), MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_10_nl
      = MUX_s_1_2_2((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_53_rtn_oreg[4]), MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_11_nl
      = MUX_s_1_2_2((MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[4]), MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_12_nl
      = MUX_s_1_2_2((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_56_rtn_oreg[4]), MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_13_nl
      = MUX_s_1_2_2((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_58_rtn_oreg[4]), MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_14_nl
      = MUX_s_1_2_2((MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_41_rtn_oreg[4]), MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_15_nl
      = MUX_s_1_2_2((MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_33_rtn_oreg[4]), MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_16_nl
      = MUX_s_1_2_2((MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_61_rtn_oreg[4]), MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_17_nl
      = MUX_s_1_2_2((MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_36_rtn_oreg[4]), MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_18_nl
      = MUX_s_1_2_2((MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_38_rtn_oreg[4]), MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_19_nl
      = MUX_s_1_2_2((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_42_rtn_oreg[4]), MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_20_nl
      = MUX_s_1_2_2((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_44_rtn_oreg[4]), MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_21_nl
      = MUX_s_1_2_2((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_46_rtn_oreg[4]), MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_22_nl
      = MUX_s_1_2_2((MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_48_rtn_oreg[4]), MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_23_nl
      = MUX_s_1_2_2((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_50_rtn_oreg[4]), MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_24_nl
      = MUX_s_1_2_2((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_52_rtn_oreg[4]), MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_25_nl
      = MUX_s_1_2_2((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_54_rtn_oreg[4]), MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_26_nl
      = MUX_s_1_2_2((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_55_rtn_oreg[4]), MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_27_nl
      = MUX_s_1_2_2((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_57_rtn_oreg[4]), MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_10_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_28_nl
      = MUX_s_1_2_2((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_59_rtn_oreg[4]), MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign MAC_1_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_nl = (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_1_sva_mx0w0!=22'b0000000000000000000000);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_qif_mux_29_nl
      = MUX_s_1_2_2((MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[0]),
      (MAC_1_leading_sign_18_1_1_0_cmp_40_rtn_oreg[4]), MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_61_nl = MUX_s_1_2_2((MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_33_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_61_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_33_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_91_nl = MUX_s_1_2_2((MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_124_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_91_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_33_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_60_nl = MUX_s_1_2_2((MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_34_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_60_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_34_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_90_nl = MUX_s_1_2_2((MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_123_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_90_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_34_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_59_nl = MUX_s_1_2_2((MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_35_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_59_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_35_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_89_nl = MUX_s_1_2_2((MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_122_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_89_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_35_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_58_nl = MUX_s_1_2_2((MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_36_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_58_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_36_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_88_nl = MUX_s_1_2_2((MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_121_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_88_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_36_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_57_nl = MUX_s_1_2_2((MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_37_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_57_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_37_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_87_nl = MUX_s_1_2_2((MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_120_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_87_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_37_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_56_nl = MUX_s_1_2_2((MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_38_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_56_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_153_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_38_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_86_nl = MUX_s_1_2_2((MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_119_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_86_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_153_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_38_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_55_nl = MUX_s_1_2_2((MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_39_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_55_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_157_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_39_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_85_nl = MUX_s_1_2_2((MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_118_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_85_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_157_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_39_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_54_nl = MUX_s_1_2_2((MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_40_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_54_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_40_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_84_nl = MUX_s_1_2_2((MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_117_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_84_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_40_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_53_nl = MUX_s_1_2_2((MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_41_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_53_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_165_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_41_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_83_nl = MUX_s_1_2_2((MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_116_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_83_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_165_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_41_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_52_nl = MUX_s_1_2_2((MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_42_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_52_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_169_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_42_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_82_nl = MUX_s_1_2_2((MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_115_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_82_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_169_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_42_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl = MUX_s_1_2_2((MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_43_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_51_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_173_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_43_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_81_nl = MUX_s_1_2_2((MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_114_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_81_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_173_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_43_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl = MUX_s_1_2_2((MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_44_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_50_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_177_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_44_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_80_nl = MUX_s_1_2_2((MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_113_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_80_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_177_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_44_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_nl = MUX_s_1_2_2((MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_45_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_49_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_181_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_45_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_79_nl = MUX_s_1_2_2((MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_112_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_79_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_181_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_45_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_48_nl = MUX_s_1_2_2((MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_46_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_48_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_185_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_46_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_78_nl = MUX_s_1_2_2((MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_111_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_78_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_185_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_46_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_47_nl = MUX_s_1_2_2((MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_47_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_47_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_189_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_47_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_77_nl = MUX_s_1_2_2((MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_110_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_77_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_189_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_47_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_46_nl = MUX_s_1_2_2((MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_48_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_46_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_193_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_48_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_76_nl = MUX_s_1_2_2((MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_109_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_76_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_193_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_48_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_45_nl = MUX_s_1_2_2((MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_49_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_45_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_197_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_49_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_75_nl = MUX_s_1_2_2((MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_108_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_75_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_197_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_49_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_44_nl = MUX_s_1_2_2((MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_50_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_44_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_201_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_50_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_74_nl = MUX_s_1_2_2((MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_107_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_74_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_201_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_50_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl = MUX_s_1_2_2((MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_51_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_43_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_205_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_51_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_73_nl = MUX_s_1_2_2((MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_106_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_73_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_205_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_51_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl = MUX_s_1_2_2((MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_52_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_42_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_209_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_52_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_72_nl = MUX_s_1_2_2((MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_105_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_72_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_209_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_52_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl = MUX_s_1_2_2((MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_53_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_41_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_213_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_53_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_71_nl = MUX_s_1_2_2((MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_104_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_71_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_213_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_53_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl = MUX_s_1_2_2((MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_54_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_40_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_217_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_54_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_70_nl = MUX_s_1_2_2((MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_103_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_70_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_217_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_54_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl = MUX_s_1_2_2((MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_55_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_39_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_221_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_55_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_69_nl = MUX_s_1_2_2((MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_102_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_69_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_221_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_55_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl = MUX_s_1_2_2((MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_56_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_38_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_225_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_56_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_68_nl = MUX_s_1_2_2((MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_101_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_68_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_225_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_56_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl = MUX_s_1_2_2((MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_57_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_37_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_229_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_57_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_67_nl = MUX_s_1_2_2((MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_100_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_67_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_229_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_57_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl = MUX_s_1_2_2((MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_58_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_36_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_233_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_58_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_66_nl = MUX_s_1_2_2((MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_99_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_66_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_233_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_58_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl = MUX_s_1_2_2((MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_59_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_35_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_237_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_59_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_65_nl = MUX_s_1_2_2((MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_98_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_65_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_237_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_59_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl = MUX_s_1_2_2((MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_60_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_34_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_241_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_60_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_64_nl = MUX_s_1_2_2((MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_97_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_64_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_241_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_60_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl = MUX_s_1_2_2((MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_61_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_33_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_245_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_61_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_63_nl = MUX_s_1_2_2((MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_96_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_63_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_245_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_61_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl = MUX_s_1_2_2((MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6]),
      (MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_62_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_32_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_249_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_62_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_62_nl = MUX_s_1_2_2((MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[5]),
      (MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_95_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_62_nl | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_249_ssc)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_62_seb;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl = MUX_v_2_2_2((MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[6:5]),
      (MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[6:5]),
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl
      = MUX_v_2_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_31_nl,
      2'b11, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_253_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_63_nl
      = MUX_v_2_2_2(2'b00, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_or_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_63_seb);
  assign and_251_nl = and_dcpl_107 & and_dcpl_225 & (~ MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_224;
  assign and_254_nl = and_dcpl_107 & and_dcpl_225 & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_224;
  assign and_257_nl = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_224;
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_63_lpi_1_dfm_6_0[3:0]);
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign and_261_nl = and_dcpl_107 & and_dcpl_235 & (~ MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_224;
  assign and_264_nl = and_dcpl_107 & and_dcpl_235 & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_224;
  assign and_267_nl = and_dcpl_107 & (~ (fsm_output[6])) & (MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_224;
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_9_lpi_1_dfm_6_0[3:0]);
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_43_nl = ~((MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_274_nl = MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_lpi_1_dfm_6_0[3:0]);
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_44_nl = ~((MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_276_nl = MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]);
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign and_279_nl = and_dcpl_108 & and_dcpl_93 & (~ (fsm_output[7])) & (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]);
  assign and_284_nl = and_dcpl_260 & and_dcpl_85 & (~((MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1));
  assign and_287_nl = and_dcpl_260 & and_dcpl_85 & (~ (MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1;
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_40_lpi_1_dfm_6_0[3:0]);
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_27_nl = ~((MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_289_nl = MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_41_lpi_1_dfm_6_0[3:0]);
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_28_nl = ~((MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_291_nl = MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_42_lpi_1_dfm_6_0[3:0]);
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_29_nl = ~((MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_293_nl = MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_43_lpi_1_dfm_6_0[3:0]);
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_30_nl = ~((MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_295_nl = MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_44_lpi_1_dfm_6_0[3:0]);
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_31_nl = ~((MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_297_nl = MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_45_lpi_1_dfm_6_0[3:0]);
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_32_nl = ~((MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_299_nl = MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_46_lpi_1_dfm_6_0[3:0]);
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_33_nl = ~((MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_301_nl = MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_47_lpi_1_dfm_6_0[3:0]);
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_34_nl = ~((MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_303_nl = MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_48_lpi_1_dfm_6_0[3:0]);
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_35_nl = ~((MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_305_nl = MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_5_lpi_1_dfm_6_0[3:0]);
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_36_nl = ~((MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_307_nl = MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_50_lpi_1_dfm_6_0[3:0]);
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_37_nl = ~((MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_309_nl = MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_51_lpi_1_dfm_6_0[3:0]);
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_39_nl = ~((MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_311_nl = MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_52_lpi_1_dfm_6_0[3:0]);
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_40_nl = ~((MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1);
  assign and_313_nl = MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_53_lpi_1_dfm_6_0[3:0]);
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_298_nl = ~(MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_315_nl = MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_54_lpi_1_dfm_6_0[3:0]);
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_299_nl = ~(MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_317_nl = MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_55_lpi_1_dfm_6_0[3:0]);
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_300_nl = ~(MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_319_nl = MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_56_lpi_1_dfm_6_0[3:0]);
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_301_nl = ~(MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_321_nl = MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_57_lpi_1_dfm_6_0[3:0]);
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_302_nl = ~(MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_323_nl = MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_58_lpi_1_dfm_6_0[3:0]);
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_303_nl = ~(MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_325_nl = MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_59_lpi_1_dfm_6_0[3:0]);
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_304_nl = ~(MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_327_nl = MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_6_lpi_1_dfm_6_0[3:0]);
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_305_nl = ~(MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_329_nl = MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_60_lpi_1_dfm_6_0[3:0]);
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_306_nl = ~(MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_331_nl = MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_61_lpi_1_dfm_6_0[3:0]);
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign nor_307_nl = ~(MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      | (MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign and_333_nl = MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_11_nl
      = MUX1HOT_s_1_67_2((MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_2_lpi_1_dfm_1_5_4[0]),
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[4]),
      (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[4]),
      (MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]), (MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[4]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[4]),
      (delay_lane_e_62_sva[4]), {and_dcpl_109 , and_573_ssc , and_575_ssc , and_579_ssc
      , and_584_ssc , and_589_ssc , and_595_ssc , and_599_ssc , and_603_ssc , and_607_ssc
      , and_613_ssc , and_617_ssc , and_621_ssc , and_625_ssc , and_631_ssc , and_635_ssc
      , and_639_ssc , and_643_ssc , and_649_ssc , and_655_ssc , and_660_ssc , and_665_ssc
      , and_669_ssc , and_673_ssc , and_677_ssc , and_681_ssc , and_685_ssc , and_689_ssc
      , and_693_ssc , and_697_ssc , and_701_ssc , and_705_ssc , and_709_ssc , and_713_ssc
      , and_718_ssc , and_722_ssc , and_726_ssc , and_730_ssc , and_735_ssc , and_739_ssc
      , and_743_ssc , and_747_ssc , and_752_ssc , and_756_ssc , and_760_ssc , and_764_ssc
      , and_769_ssc , and_773_ssc , and_777_ssc , and_781_ssc , and_785_ssc , and_789_ssc
      , and_793_ssc , and_797_ssc , and_801_ssc , and_805_ssc , and_809_ssc , and_813_ssc
      , and_817_ssc , and_821_ssc , and_825_ssc , and_829_ssc , and_833_ssc , and_837_ssc
      , and_841_ssc , and_845_ssc , and_dcpl_207});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_and_nl
      = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_11_nl
      & (~ and_568_ssc);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl
      = MUX_v_4_2_2(4'b0000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_33_nl
      = MUX1HOT_v_4_67_2((MAC_1_leading_sign_18_1_1_0_cmp_63_rtn_oreg[3:0]), ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_126_nl,
      MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1, (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_10_sva_rsp_2[3:0]),
      (MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_34_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_56_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[3:0]),
      (MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_1_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]), (MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]), (MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_34_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_35_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_36_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_37_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_38_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_39_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]), (MAC_40_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_35_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_36_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_37_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_38_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_39_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_58_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_59_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0[3:0]),
      (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_lpi_1_dfm_4_0[3:0]),
      (delay_lane_e_62_sva[3:0]), {and_dcpl_109 , and_573_ssc , and_575_ssc , and_579_ssc
      , and_584_ssc , and_589_ssc , and_595_ssc , and_599_ssc , and_603_ssc , and_607_ssc
      , and_613_ssc , and_617_ssc , and_621_ssc , and_625_ssc , and_631_ssc , and_635_ssc
      , and_639_ssc , and_643_ssc , and_649_ssc , and_655_ssc , and_660_ssc , and_665_ssc
      , and_669_ssc , and_673_ssc , and_677_ssc , and_681_ssc , and_685_ssc , and_689_ssc
      , and_693_ssc , and_697_ssc , and_701_ssc , and_705_ssc , and_709_ssc , and_713_ssc
      , and_718_ssc , and_722_ssc , and_726_ssc , and_730_ssc , and_735_ssc , and_739_ssc
      , and_743_ssc , and_747_ssc , and_752_ssc , and_756_ssc , and_760_ssc , and_764_ssc
      , and_769_ssc , and_773_ssc , and_777_ssc , and_781_ssc , and_785_ssc , and_789_ssc
      , and_793_ssc , and_797_ssc , and_801_ssc , and_805_ssc , and_809_ssc , and_813_ssc
      , and_817_ssc , and_821_ssc , and_825_ssc , and_829_ssc , and_833_ssc , and_837_ssc
      , and_841_ssc , and_845_ssc , and_dcpl_207});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_or_nl
      = MUX_v_4_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_1_mux1h_33_nl,
      4'b1111, and_568_ssc);
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_1_nl = or_770_rgt & and_118_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_4_nl = or_756_rgt & and_119_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_7_nl = or_749_rgt & and_120_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_10_nl = or_743_rgt & and_121_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_13_nl = or_737_rgt & and_122_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_16_nl = or_729_rgt & nor_248_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_19_nl = or_723_rgt & and_125_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_22_nl = or_717_rgt & and_127_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_25_nl = or_710_rgt & and_129_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_28_nl = or_704_rgt & and_133_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_31_nl = or_697_rgt & and_135_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_34_nl = or_683_rgt & and_137_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_37_nl = or_675_rgt & and_138_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_40_nl = or_667_rgt & and_139_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_43_nl = or_660_rgt & and_140_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_46_nl = or_653_rgt & and_141_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_49_nl = or_646_rgt & and_142_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_52_nl = or_639_rgt & and_143_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_55_nl = or_631_rgt & and_144_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_58_nl = or_470_rgt & and_145_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_61_nl = or_453_rgt & and_146_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_64_nl = or_445_rgt & and_149_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_67_nl = or_437_rgt & and_151_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_70_nl = or_430_rgt & and_153_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_73_nl = or_422_rgt & and_155_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_76_nl = or_415_rgt & and_156_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_79_nl = or_408_rgt & and_158_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_82_nl = or_401_rgt & and_159_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_85_nl = or_763_rgt & and_160_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_88_nl = or_690_rgt & and_161_rgt;
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_and_91_nl = or_462_rgt & and_162_rgt;
  assign MAC_10_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_nl
      = ~((ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva_mx0w0[3:0]!=4'b0000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_nl = (~
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      & and_dcpl_109;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_and_1_nl =
      MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & and_dcpl_109;
  assign and_1933_nl = (fsm_output[7]) & (~((MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp));
  assign nand_88_nl = ~((MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_89_nl = ~((MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1103_nl = MUX_s_1_2_2(nand_88_nl, nand_89_nl, fsm_output[7]);
  assign mux_1104_nl = MUX_s_1_2_2(and_1933_nl, mux_1103_nl, fsm_output[6]);
  assign nand_90_nl = ~((MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_91_nl = ~((MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1101_nl = MUX_s_1_2_2(nand_90_nl, nand_91_nl, fsm_output[7]);
  assign nand_92_nl = ~((MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_93_nl = ~((MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1100_nl = MUX_s_1_2_2(nand_92_nl, nand_93_nl, fsm_output[7]);
  assign mux_1102_nl = MUX_s_1_2_2(mux_1101_nl, mux_1100_nl, fsm_output[6]);
  assign mux_1105_nl = MUX_s_1_2_2(mux_1104_nl, mux_1102_nl, fsm_output[2]);
  assign nand_94_nl = ~((MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_95_nl = ~((MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1097_nl = MUX_s_1_2_2(nand_94_nl, nand_95_nl, fsm_output[7]);
  assign nand_96_nl = ~((MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_97_nl = ~((MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1096_nl = MUX_s_1_2_2(nand_96_nl, nand_97_nl, fsm_output[7]);
  assign mux_1098_nl = MUX_s_1_2_2(mux_1097_nl, mux_1096_nl, fsm_output[6]);
  assign nand_98_nl = ~((MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_99_nl = ~((MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1094_nl = MUX_s_1_2_2(nand_98_nl, nand_99_nl, fsm_output[7]);
  assign nand_100_nl = ~((MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_101_nl = ~((MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1093_nl = MUX_s_1_2_2(nand_100_nl, nand_101_nl, fsm_output[7]);
  assign mux_1095_nl = MUX_s_1_2_2(mux_1094_nl, mux_1093_nl, fsm_output[6]);
  assign mux_1099_nl = MUX_s_1_2_2(mux_1098_nl, mux_1095_nl, fsm_output[2]);
  assign mux_1106_nl = MUX_s_1_2_2(mux_1105_nl, mux_1099_nl, fsm_output[3]);
  assign nand_102_nl = ~((MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_103_nl = ~((MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1089_nl = MUX_s_1_2_2(nand_102_nl, nand_103_nl, fsm_output[7]);
  assign nand_104_nl = ~((MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_105_nl = ~((MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1088_nl = MUX_s_1_2_2(nand_104_nl, nand_105_nl, fsm_output[7]);
  assign mux_1090_nl = MUX_s_1_2_2(mux_1089_nl, mux_1088_nl, fsm_output[6]);
  assign nand_106_nl = ~((MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_107_nl = ~((MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1086_nl = MUX_s_1_2_2(nand_106_nl, nand_107_nl, fsm_output[7]);
  assign nand_108_nl = ~((MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_109_nl = ~((MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1085_nl = MUX_s_1_2_2(nand_108_nl, nand_109_nl, fsm_output[7]);
  assign mux_1087_nl = MUX_s_1_2_2(mux_1086_nl, mux_1085_nl, fsm_output[6]);
  assign mux_1091_nl = MUX_s_1_2_2(mux_1090_nl, mux_1087_nl, fsm_output[2]);
  assign nand_110_nl = ~((MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_111_nl = ~((MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1082_nl = MUX_s_1_2_2(nand_110_nl, nand_111_nl, fsm_output[7]);
  assign nand_112_nl = ~((MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_113_nl = ~((MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1081_nl = MUX_s_1_2_2(nand_112_nl, nand_113_nl, fsm_output[7]);
  assign mux_1083_nl = MUX_s_1_2_2(mux_1082_nl, mux_1081_nl, fsm_output[6]);
  assign nand_114_nl = ~((MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_115_nl = ~((MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1079_nl = MUX_s_1_2_2(nand_114_nl, nand_115_nl, fsm_output[7]);
  assign nand_116_nl = ~((MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_117_nl = ~((MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1078_nl = MUX_s_1_2_2(nand_116_nl, nand_117_nl, fsm_output[7]);
  assign mux_1080_nl = MUX_s_1_2_2(mux_1079_nl, mux_1078_nl, fsm_output[6]);
  assign mux_1084_nl = MUX_s_1_2_2(mux_1083_nl, mux_1080_nl, fsm_output[2]);
  assign mux_1092_nl = MUX_s_1_2_2(mux_1091_nl, mux_1084_nl, fsm_output[3]);
  assign mux_1107_nl = MUX_s_1_2_2(mux_1106_nl, mux_1092_nl, fsm_output[4]);
  assign nand_118_nl = ~((MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_119_nl = ~((MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1073_nl = MUX_s_1_2_2(nand_118_nl, nand_119_nl, fsm_output[7]);
  assign nand_120_nl = ~((MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_121_nl = ~((MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1072_nl = MUX_s_1_2_2(nand_120_nl, nand_121_nl, fsm_output[7]);
  assign mux_1074_nl = MUX_s_1_2_2(mux_1073_nl, mux_1072_nl, fsm_output[6]);
  assign nand_122_nl = ~((MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_123_nl = ~((MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1070_nl = MUX_s_1_2_2(nand_122_nl, nand_123_nl, fsm_output[7]);
  assign nand_124_nl = ~((MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_125_nl = ~((MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1069_nl = MUX_s_1_2_2(nand_124_nl, nand_125_nl, fsm_output[7]);
  assign mux_1071_nl = MUX_s_1_2_2(mux_1070_nl, mux_1069_nl, fsm_output[6]);
  assign mux_1075_nl = MUX_s_1_2_2(mux_1074_nl, mux_1071_nl, fsm_output[2]);
  assign nand_126_nl = ~((MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_127_nl = ~((MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1066_nl = MUX_s_1_2_2(nand_126_nl, nand_127_nl, fsm_output[7]);
  assign nand_128_nl = ~((MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_129_nl = ~((MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1065_nl = MUX_s_1_2_2(nand_128_nl, nand_129_nl, fsm_output[7]);
  assign mux_1067_nl = MUX_s_1_2_2(mux_1066_nl, mux_1065_nl, fsm_output[6]);
  assign nand_130_nl = ~((MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_131_nl = ~((MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1063_nl = MUX_s_1_2_2(nand_130_nl, nand_131_nl, fsm_output[7]);
  assign nand_132_nl = ~((MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_133_nl = ~((MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1062_nl = MUX_s_1_2_2(nand_132_nl, nand_133_nl, fsm_output[7]);
  assign mux_1064_nl = MUX_s_1_2_2(mux_1063_nl, mux_1062_nl, fsm_output[6]);
  assign mux_1068_nl = MUX_s_1_2_2(mux_1067_nl, mux_1064_nl, fsm_output[2]);
  assign mux_1076_nl = MUX_s_1_2_2(mux_1075_nl, mux_1068_nl, fsm_output[3]);
  assign nand_134_nl = ~((MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_135_nl = ~((MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1058_nl = MUX_s_1_2_2(nand_134_nl, nand_135_nl, fsm_output[7]);
  assign nand_136_nl = ~((MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_137_nl = ~((MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1057_nl = MUX_s_1_2_2(nand_136_nl, nand_137_nl, fsm_output[7]);
  assign mux_1059_nl = MUX_s_1_2_2(mux_1058_nl, mux_1057_nl, fsm_output[6]);
  assign nand_138_nl = ~((MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_139_nl = ~((MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1055_nl = MUX_s_1_2_2(nand_138_nl, nand_139_nl, fsm_output[7]);
  assign nand_140_nl = ~((MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_141_nl = ~((MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1054_nl = MUX_s_1_2_2(nand_140_nl, nand_141_nl, fsm_output[7]);
  assign mux_1056_nl = MUX_s_1_2_2(mux_1055_nl, mux_1054_nl, fsm_output[6]);
  assign mux_1060_nl = MUX_s_1_2_2(mux_1059_nl, mux_1056_nl, fsm_output[2]);
  assign nand_142_nl = ~((MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_143_nl = ~((MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1051_nl = MUX_s_1_2_2(nand_142_nl, nand_143_nl, fsm_output[7]);
  assign nand_144_nl = ~((MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_145_nl = ~((MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1050_nl = MUX_s_1_2_2(nand_144_nl, nand_145_nl, fsm_output[7]);
  assign mux_1052_nl = MUX_s_1_2_2(mux_1051_nl, mux_1050_nl, fsm_output[6]);
  assign nand_146_nl = ~((MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_147_nl = ~((MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1048_nl = MUX_s_1_2_2(nand_146_nl, nand_147_nl, fsm_output[7]);
  assign nand_148_nl = ~((MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign nand_149_nl = ~((MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp);
  assign mux_1047_nl = MUX_s_1_2_2(nand_148_nl, nand_149_nl, fsm_output[7]);
  assign mux_1049_nl = MUX_s_1_2_2(mux_1048_nl, mux_1047_nl, fsm_output[6]);
  assign mux_1053_nl = MUX_s_1_2_2(mux_1052_nl, mux_1049_nl, fsm_output[2]);
  assign mux_1061_nl = MUX_s_1_2_2(mux_1060_nl, mux_1053_nl, fsm_output[3]);
  assign mux_1077_nl = MUX_s_1_2_2(mux_1076_nl, mux_1061_nl, fsm_output[4]);
  assign mux_1108_nl = MUX_s_1_2_2(mux_1107_nl, mux_1077_nl, fsm_output[5]);
  assign nand_150_nl = ~((fsm_output[1]) & mux_1108_nl);
  assign nor_845_nl = ~((fsm_output[7:2]!=6'b000000));
  assign mux_1109_nl = MUX_s_1_2_2(nand_150_nl, nor_845_nl, fsm_output[0]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_33_nl
      = ~((~ MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_66_nl
      = MUX1HOT_v_5_3_2((MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_34_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_33_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_133_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_94_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_66_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_33_seb);
  assign nor_640_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm
      | (~ and_1698_cse));
  assign or_1036_nl = nor_641_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[6]);
  assign mux_655_nl = MUX_s_1_2_2(nor_640_nl, and_1698_cse, or_1036_nl);
  assign nor_642_nl = ~((fsm_output[2]) | mux_655_nl);
  assign mux_656_nl = MUX_s_1_2_2(nor_642_nl, nor_tmp, fsm_output[3]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_312_nl = (mux_656_nl
      | or_dcpl_278) & and_184_ssc;
  assign and_1301_nl = ((~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_itm)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_6_tmp[6])
      | nor_641_cse) & and_dcpl_497 & and_184_ssc;
  assign mux_657_nl = MUX_s_1_2_2((fsm_output[2]), (~ nor_tmp), fsm_output[3]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_34_nl
      = ~((~ MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_68_nl
      = MUX1HOT_v_5_3_2((MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_35_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_34_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_137_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_93_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_68_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_34_seb);
  assign or_995_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6
      | nor_616_cse | (fsm_output[7]);
  assign mux_636_nl = MUX_s_1_2_2((fsm_output[7]), or_995_nl, and_1698_cse);
  assign nor_617_nl = ~((fsm_output[4:3]!=2'b00) | mux_636_nl);
  assign and_1733_nl = (fsm_output[3]) & (fsm_output[4]) & (fsm_output[1]) & (fsm_output[7]);
  assign mux_637_nl = MUX_s_1_2_2(nor_617_nl, and_1733_nl, fsm_output[2]);
  assign or_991_nl = (fsm_output[6:5]!=2'b00);
  assign mux_638_nl = MUX_s_1_2_2(mux_637_nl, (fsm_output[7]), or_991_nl);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_310_nl = (mux_638_nl
      | (fsm_output[8])) & nor_252_ssc;
  assign and_1277_nl = and_dcpl_497 & (nor_616_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_40_lpi_1_dfm_6)
      & nor_252_ssc;
  assign mux_639_nl = MUX_s_1_2_2(not_tmp_640, or_tmp_227, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_35_nl
      = ~((~ MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_70_nl
      = MUX1HOT_v_5_3_2((MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_36_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_35_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_141_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_92_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_70_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_35_seb);
  assign nor_612_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_633_nl = MUX_s_1_2_2(nor_612_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6);
  assign nor_613_nl = ~((fsm_output[6:2]!=5'b00000) | mux_633_nl);
  assign mux_634_nl = MUX_s_1_2_2(nor_613_nl, mux_tmp_213, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_308_nl = (mux_634_nl
      | (fsm_output[8])) & nor_253_ssc;
  assign and_1273_nl = (nor_614_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_41_lpi_1_dfm_6)
      & and_dcpl_497 & nor_253_ssc;
  assign mux_635_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_213, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_36_nl
      = ~((~ MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_72_nl
      = MUX1HOT_v_5_3_2((MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_37_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_36_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_145_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_91_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_72_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_36_seb);
  assign nor_608_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_630_nl = MUX_s_1_2_2(nor_608_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6);
  assign nor_609_nl = ~((fsm_output[6:2]!=5'b00000) | mux_630_nl);
  assign mux_631_nl = MUX_s_1_2_2(nor_609_nl, mux_tmp_215, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_306_nl = (mux_631_nl
      | (fsm_output[8])) & nor_254_ssc;
  assign and_1269_nl = (nor_610_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_42_lpi_1_dfm_6)
      & and_dcpl_497 & nor_254_ssc;
  assign mux_632_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_215, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_37_nl
      = ~((~ MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_74_nl
      = MUX1HOT_v_5_3_2((MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_38_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_37_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_149_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_90_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_74_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_37_seb);
  assign nor_604_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
      | (~ and_1698_cse));
  assign mux_627_nl = MUX_s_1_2_2(nor_604_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6);
  assign nor_605_nl = ~((fsm_output[6:2]!=5'b00000) | mux_627_nl);
  assign mux_628_nl = MUX_s_1_2_2(nor_605_nl, mux_tmp_217, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_304_nl = (mux_628_nl
      | (fsm_output[8])) & nor_255_ssc;
  assign and_1265_nl = (nor_606_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_6)
      & and_dcpl_497 & nor_255_ssc;
  assign mux_629_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_217, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_38_nl
      = ~((~ MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_76_nl
      = MUX1HOT_v_5_3_2((MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_39_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_38_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_153_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_89_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_76_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_38_seb);
  assign or_968_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6
      | nor_600_cse | (fsm_output[5]) | (fsm_output[7]);
  assign mux_622_nl = MUX_s_1_2_2(or_969_cse, or_968_nl, and_1698_cse);
  assign nor_601_nl = ~((fsm_output[3]) | mux_622_nl);
  assign and_1730_nl = (fsm_output[3]) & (fsm_output[1]) & (fsm_output[5]) & (fsm_output[7]);
  assign mux_623_nl = MUX_s_1_2_2(nor_601_nl, and_1730_nl, fsm_output[2]);
  assign mux_624_nl = MUX_s_1_2_2(mux_623_nl, and_1731_cse, fsm_output[4]);
  assign mux_625_nl = MUX_s_1_2_2(mux_624_nl, (fsm_output[7]), fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_302_nl = (mux_625_nl
      | (fsm_output[8])) & nor_256_ssc;
  assign and_1261_nl = and_dcpl_497 & (nor_600_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_44_lpi_1_dfm_6)
      & nor_256_ssc;
  assign mux_626_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_219, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_39_nl
      = ~((~ MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_78_nl
      = MUX1HOT_v_5_3_2((MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_39_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_157_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_88_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_78_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_39_seb);
  assign nor_596_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_619_nl = MUX_s_1_2_2(nor_596_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6);
  assign nor_597_nl = ~((fsm_output[6:2]!=5'b00000) | mux_619_nl);
  assign mux_620_nl = MUX_s_1_2_2(nor_597_nl, mux_tmp_221, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_300_nl = (mux_620_nl
      | (fsm_output[8])) & nor_257_ssc;
  assign and_1257_nl = (nor_598_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_45_lpi_1_dfm_6)
      & and_dcpl_497 & nor_257_ssc;
  assign mux_621_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_221, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_40_nl
      = ~((~ MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_80_nl
      = MUX1HOT_v_5_3_2((MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_41_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_40_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_161_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_87_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_80_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_40_seb);
  assign nor_592_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_5
      | (~ and_1698_cse));
  assign mux_616_nl = MUX_s_1_2_2(nor_592_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6);
  assign nor_593_nl = ~((fsm_output[6:2]!=5'b00000) | mux_616_nl);
  assign mux_617_nl = MUX_s_1_2_2(nor_593_nl, mux_tmp_223, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_298_nl = (mux_617_nl
      | (fsm_output[8])) & nor_258_ssc;
  assign and_1253_nl = (nor_594_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_46_lpi_1_dfm_6)
      & and_dcpl_497 & nor_258_ssc;
  assign mux_618_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_223, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_41_nl
      = ~((~ MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_82_nl
      = MUX1HOT_v_5_3_2((MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_42_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_41_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_165_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_86_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_82_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_41_seb);
  assign or_950_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6
      | nor_587_cse | (fsm_output[7]);
  assign mux_612_nl = MUX_s_1_2_2((fsm_output[7]), or_950_nl, and_1698_cse);
  assign nor_588_nl = ~((fsm_output[4]) | (fsm_output[5]) | (fsm_output[2]) | mux_612_nl);
  assign and_1246_nl = (fsm_output[5:4]==2'b11) & or_1164_cse & (fsm_output[7]);
  assign mux_613_nl = MUX_s_1_2_2(nor_588_nl, and_1246_nl, fsm_output[3]);
  assign mux_614_nl = MUX_s_1_2_2(mux_613_nl, (fsm_output[7]), fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_296_nl = (mux_614_nl
      | (fsm_output[8])) & nor_259_ssc;
  assign and_1249_nl = and_dcpl_497 & (nor_587_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_47_lpi_1_dfm_6)
      & nor_259_ssc;
  assign mux_615_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_225, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_42_nl
      = ~((~ MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_84_nl
      = MUX1HOT_v_5_3_2((MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_43_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_42_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_169_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_85_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_84_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_42_seb);
  assign nor_583_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_5
      | (~ and_1698_cse));
  assign mux_609_nl = MUX_s_1_2_2(nor_583_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6);
  assign nor_584_nl = ~((fsm_output[6:2]!=5'b00000) | mux_609_nl);
  assign mux_610_nl = MUX_s_1_2_2(nor_584_nl, mux_tmp_227, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_294_nl = (mux_610_nl
      | (fsm_output[8])) & nor_260_ssc;
  assign and_1244_nl = (nor_585_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_48_lpi_1_dfm_6)
      & and_dcpl_497 & nor_260_ssc;
  assign mux_611_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_227, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_43_nl
      = ~((~ MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_86_nl
      = MUX1HOT_v_5_3_2((MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_44_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_43_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_173_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_84_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_86_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_43_seb);
  assign or_935_nl = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_4_0[4])
      | (~ (fsm_output[1])))) | (fsm_output[5:2]!=4'b0000);
  assign mux_605_nl = MUX_s_1_2_2(or_935_nl, or_tmp_589, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6);
  assign mux_606_nl = MUX_s_1_2_2(or_456_cse, mux_605_nl, fsm_output[0]);
  assign nor_580_nl = ~((fsm_output[7]) | mux_606_nl);
  assign and_1237_nl = (fsm_output[7]) & or_tmp_589;
  assign mux_607_nl = MUX_s_1_2_2(nor_580_nl, and_1237_nl, fsm_output[6]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_292_nl = (mux_607_nl
      | (fsm_output[8])) & nor_261_ssc;
  assign and_1240_nl = and_dcpl_497 & (nor_581_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_49_lpi_1_dfm_6)
      & nor_261_ssc;
  assign mux_608_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_229, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_44_nl
      = ~((~ MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_88_nl
      = MUX1HOT_v_5_3_2((MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_45_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_44_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_177_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_83_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_88_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_44_seb);
  assign and_1738_nl = (nor_636_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[6]))
      & (fsm_output[1:0]==2'b11);
  assign mux_652_nl = MUX_s_1_2_2(and_1698_cse, and_1738_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm);
  assign nor_638_nl = ~((fsm_output[3:2]!=2'b00) | mux_652_nl);
  assign mux_653_nl = MUX_s_1_2_2(nor_638_nl, or_dcpl_115, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_291_nl = (mux_653_nl
      | or_dcpl_368) & and_196_ssc;
  assign and_1297_nl = (nor_636_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_8_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_itm))
      & and_dcpl_497 & and_196_ssc;
  assign mux_654_nl = MUX_s_1_2_2(nor_136_cse, or_dcpl_115, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_45_nl
      = ~((~ MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_90_nl
      = MUX1HOT_v_5_3_2((MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_46_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_45_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_181_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_82_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_90_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_45_seb);
  assign nor_576_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_602_nl = MUX_s_1_2_2(nor_576_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6);
  assign nor_577_nl = ~((fsm_output[6:2]!=5'b00000) | mux_602_nl);
  assign mux_603_nl = MUX_s_1_2_2(nor_577_nl, mux_tmp_232, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_289_nl = (mux_603_nl
      | (fsm_output[8])) & nor_262_ssc;
  assign and_1235_nl = (nor_578_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_50_lpi_1_dfm_6)
      & and_dcpl_497 & nor_262_ssc;
  assign mux_604_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_232, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_46_nl
      = ~((~ MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_92_nl
      = MUX1HOT_v_5_3_2((MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_47_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_46_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_185_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_81_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_92_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_46_seb);
  assign nor_572_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_599_nl = MUX_s_1_2_2(nor_572_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6);
  assign nor_573_nl = ~((fsm_output[6:2]!=5'b00000) | mux_599_nl);
  assign mux_600_nl = MUX_s_1_2_2(nor_573_nl, mux_tmp_234, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_287_nl = (mux_600_nl
      | (fsm_output[8])) & nor_263_ssc;
  assign and_1231_nl = (nor_574_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_51_lpi_1_dfm_6)
      & and_dcpl_497 & nor_263_ssc;
  assign mux_601_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_234, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_nl
      = ~((~ MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_94_nl
      = MUX1HOT_v_5_3_2((MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_48_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_47_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_189_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_80_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_94_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_47_seb);
  assign or_917_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6
      | nor_568_cse | (fsm_output[7:6]!=2'b00);
  assign mux_595_nl = MUX_s_1_2_2(or_918_cse, or_917_nl, and_1698_cse);
  assign nor_569_nl = ~((fsm_output[3]) | mux_595_nl);
  assign and_1724_nl = (fsm_output[3]) & (fsm_output[1]) & (fsm_output[6]) & (fsm_output[7]);
  assign mux_596_nl = MUX_s_1_2_2(nor_569_nl, and_1724_nl, fsm_output[2]);
  assign mux_597_nl = MUX_s_1_2_2(mux_596_nl, and_1725_cse, or_627_cse);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_285_nl = (mux_597_nl
      | (fsm_output[8])) & nor_264_ssc;
  assign and_1227_nl = and_dcpl_497 & (nor_568_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_52_lpi_1_dfm_6)
      & nor_264_ssc;
  assign mux_598_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_236, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_48_nl
      = ~((~ MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_96_nl
      = MUX1HOT_v_5_3_2((MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_49_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_48_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_193_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_79_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_96_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_48_seb);
  assign nor_564_nl = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_4_0[4])
      | (~ and_1698_cse));
  assign mux_592_nl = MUX_s_1_2_2(nor_564_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6);
  assign nor_565_nl = ~((fsm_output[6:2]!=5'b00000) | mux_592_nl);
  assign mux_593_nl = MUX_s_1_2_2(nor_565_nl, mux_tmp_238, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_283_nl = (mux_593_nl
      | (fsm_output[8])) & nor_265_ssc;
  assign and_1223_nl = (nor_566_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_53_lpi_1_dfm_6)
      & and_dcpl_497 & nor_265_ssc;
  assign mux_594_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_238, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_49_nl
      = ~((~ MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_98_nl
      = MUX1HOT_v_5_3_2((MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_50_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_49_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_197_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_78_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_98_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_49_seb);
  assign nor_560_nl = ~((ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0[4])
      | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
      | (~ and_1698_cse));
  assign mux_589_nl = MUX_s_1_2_2(nor_560_nl, and_1698_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6);
  assign nor_561_nl = ~((fsm_output[6:2]!=5'b00000) | mux_589_nl);
  assign mux_590_nl = MUX_s_1_2_2(nor_561_nl, mux_tmp_240, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_281_nl = (mux_590_nl
      | (fsm_output[8])) & nor_266_ssc;
  assign and_1219_nl = (nor_562_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_6)
      & and_dcpl_497 & nor_266_ssc;
  assign mux_591_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_240, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_50_nl
      = ~((~ MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_100_nl
      = MUX1HOT_v_5_3_2((MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_51_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_50_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_201_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_77_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_100_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_50_seb);
  assign or_897_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6
      | nor_555_cse | (fsm_output[7:6]!=2'b00);
  assign mux_585_nl = MUX_s_1_2_2(or_918_cse, or_897_nl, and_1698_cse);
  assign nor_556_nl = ~((fsm_output[4]) | (fsm_output[2]) | mux_585_nl);
  assign and_1212_nl = (fsm_output[4]) & or_1164_cse & (fsm_output[7:6]==2'b11);
  assign mux_586_nl = MUX_s_1_2_2(nor_556_nl, and_1212_nl, fsm_output[3]);
  assign mux_587_nl = MUX_s_1_2_2(mux_586_nl, and_1725_cse, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_279_nl = (mux_587_nl
      | (fsm_output[8])) & nor_267_ssc;
  assign and_1215_nl = and_dcpl_497 & (nor_555_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_55_lpi_1_dfm_6)
      & nor_267_ssc;
  assign mux_588_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_242, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_51_nl
      = ~((~ MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_102_nl
      = MUX1HOT_v_5_3_2((MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_52_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_51_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_205_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_76_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_102_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_51_seb);
  assign nor_552_nl = ~((fsm_output[6:2]!=5'b00000) | (or_1162_cse & (fsm_output[1:0]==2'b11)));
  assign mux_583_nl = MUX_s_1_2_2(nor_552_nl, mux_tmp_244, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_277_nl = (mux_583_nl
      | (fsm_output[8])) & nor_268_ssc;
  assign and_1210_nl = or_1162_cse & and_dcpl_497 & nor_268_ssc;
  assign mux_584_nl = MUX_s_1_2_2(not_tmp_640, mux_tmp_244, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_52_nl
      = ~((~ MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_104_nl
      = MUX1HOT_v_5_3_2((MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_53_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_52_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_209_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_75_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_104_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_52_seb);
  assign or_882_nl = (~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_4_0[4])
      | (~ (fsm_output[1])))) | (fsm_output[4:2]!=3'b000);
  assign mux_579_nl = MUX_s_1_2_2(or_882_nl, or_1113_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6);
  assign mux_580_nl = MUX_s_1_2_2(or_452_cse, mux_579_nl, fsm_output[0]);
  assign nor_547_nl = ~((fsm_output[7:6]!=2'b00) | mux_580_nl);
  assign and_1203_nl = (fsm_output[7:6]==2'b11) & or_1113_cse;
  assign mux_581_nl = MUX_s_1_2_2(nor_547_nl, and_1203_nl, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_275_nl = (mux_581_nl
      | (fsm_output[8])) & nor_269_ssc;
  assign and_1206_nl = (nor_548_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_57_lpi_1_dfm_6)
      & and_dcpl_497 & nor_269_ssc;
  assign mux_582_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_16, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_53_nl
      = ~((~ MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_106_nl
      = MUX1HOT_v_5_3_2((MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_54_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_53_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_213_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_74_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_106_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_53_seb);
  assign nor_544_nl = ~((fsm_output[6:2]!=5'b00000) | (or_1161_cse & (fsm_output[1:0]==2'b11)));
  assign mux_577_nl = MUX_s_1_2_2(nor_544_nl, and_tmp_17, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_273_nl = (mux_577_nl
      | (fsm_output[8])) & nor_270_ssc;
  assign and_1201_nl = or_1161_cse & and_dcpl_497 & nor_270_ssc;
  assign mux_578_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_17, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_54_nl
      = ~((~ MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_108_nl
      = MUX1HOT_v_5_3_2((MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_55_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_54_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_217_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_73_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_108_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_54_seb);
  assign nor_539_nl = ~((fsm_output[6:2]!=5'b00000) | (or_1160_cse & (fsm_output[1:0]==2'b11)));
  assign mux_575_nl = MUX_s_1_2_2(nor_539_nl, and_tmp_18, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_271_nl = (mux_575_nl
      | (fsm_output[8])) & nor_271_ssc;
  assign and_1197_nl = or_1160_cse & and_dcpl_497 & nor_271_ssc;
  assign mux_576_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_18, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_55_nl
      = ~((~ MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_110_nl
      = MUX1HOT_v_5_3_2((MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_56_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_55_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_221_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_72_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_110_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_55_seb);
  assign and_1737_nl = (nor_632_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[6]))
      & (fsm_output[1:0]==2'b11);
  assign mux_649_nl = MUX_s_1_2_2(and_1698_cse, and_1737_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm);
  assign nor_634_nl = ~((fsm_output[3:2]!=2'b00) | mux_649_nl);
  assign mux_650_nl = MUX_s_1_2_2(nor_634_nl, or_123_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_270_nl = (mux_650_nl
      | or_dcpl_368) & and_210_ssc;
  assign and_1293_nl = (nor_632_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_10_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_itm))
      & and_dcpl_497 & and_210_ssc;
  assign mux_651_nl = MUX_s_1_2_2(nor_136_cse, or_123_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_56_nl
      = ~((~ MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_112_nl
      = MUX1HOT_v_5_3_2((MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_57_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_56_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_225_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_71_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_112_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_56_seb);
  assign or_864_nl = (fsm_output[7:5]!=3'b000);
  assign or_863_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6
      | nor_533_cse | (fsm_output[7:5]!=3'b000);
  assign mux_571_nl = MUX_s_1_2_2(or_864_nl, or_863_nl, and_1698_cse);
  assign nor_534_nl = ~((fsm_output[3]) | mux_571_nl);
  assign and_1714_nl = (fsm_output[3]) & (fsm_output[1]) & (fsm_output[5]) & (fsm_output[6])
      & (fsm_output[7]);
  assign mux_572_nl = MUX_s_1_2_2(nor_534_nl, and_1714_nl, fsm_output[2]);
  assign and_1715_nl = (fsm_output[7:5]==3'b111);
  assign mux_573_nl = MUX_s_1_2_2(mux_572_nl, and_1715_nl, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_268_nl = (mux_573_nl
      | (fsm_output[8])) & nor_272_ssc;
  assign and_1193_nl = (nor_533_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_6)
      & and_dcpl_497 & nor_272_ssc;
  assign mux_574_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_19, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_57_nl
      = ~((~ MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_114_nl
      = MUX1HOT_v_5_3_2((MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_58_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_57_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_229_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_70_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_114_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_57_seb);
  assign nor_530_nl = ~((fsm_output[6:2]!=5'b00000) | (or_1159_cse & (fsm_output[1:0]==2'b11)));
  assign mux_569_nl = MUX_s_1_2_2(nor_530_nl, and_tmp_20, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_266_nl = (mux_569_nl
      | (fsm_output[8])) & nor_273_ssc;
  assign and_1189_nl = or_1159_cse & and_dcpl_497 & nor_273_ssc;
  assign mux_570_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_20, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_58_nl
      = ~((~ MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_116_nl
      = MUX1HOT_v_5_3_2((MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_59_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_58_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_233_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_69_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_116_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_58_seb);
  assign nor_525_nl = ~((fsm_output[6:2]!=5'b00000) | (or_1158_cse & (fsm_output[1:0]==2'b11)));
  assign mux_567_nl = MUX_s_1_2_2(nor_525_nl, and_tmp_21, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_264_nl = (mux_567_nl
      | (fsm_output[8])) & nor_274_ssc;
  assign and_1185_nl = or_1158_cse & and_dcpl_497 & nor_274_ssc;
  assign mux_568_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_21, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_59_nl
      = ~((~ MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_118_nl
      = MUX1HOT_v_5_3_2((MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_60_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_59_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_237_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_68_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_118_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_59_seb);
  assign nor_520_nl = ~((fsm_output[7:3]!=5'b00000));
  assign or_844_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0[4]);
  assign mux_561_nl = MUX_s_1_2_2(and_1695_cse, mux_tmp_557, or_844_nl);
  assign mux_562_nl = MUX_s_1_2_2(mux_561_nl, and_1695_cse, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6);
  assign mux_563_nl = MUX_s_1_2_2(mux_tmp_557, mux_562_nl, fsm_output[0]);
  assign mux_564_nl = MUX_s_1_2_2(nor_520_nl, mux_563_nl, fsm_output[1]);
  assign mux_565_nl = MUX_s_1_2_2(mux_564_nl, and_1695_cse, fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_262_nl = (mux_565_nl
      | (fsm_output[8])) & nor_275_ssc;
  assign and_1181_nl = (nor_521_cse | ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_6)
      & and_dcpl_497 & nor_275_ssc;
  assign mux_566_nl = MUX_s_1_2_2(not_tmp_640, and_tmp_22, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_60_nl
      = ~((~ MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_120_nl
      = MUX1HOT_v_5_3_2((MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_61_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_60_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_241_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_67_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_120_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_60_seb);
  assign and_1736_nl = (nor_628_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[6]))
      & (fsm_output[1:0]==2'b11);
  assign mux_646_nl = MUX_s_1_2_2(and_1698_cse, and_1736_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm);
  assign nor_630_nl = ~((fsm_output[3:2]!=2'b00) | mux_646_nl);
  assign mux_647_nl = MUX_s_1_2_2(nor_630_nl, and_4_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_261_nl = (mux_647_nl
      | or_dcpl_368) & and_219_ssc;
  assign and_1289_nl = (nor_628_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_12_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_itm))
      & and_dcpl_497 & and_219_ssc;
  assign mux_648_nl = MUX_s_1_2_2(nor_136_cse, and_4_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_61_nl
      = ~((~ MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_122_nl
      = MUX1HOT_v_5_3_2((MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_62_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_61_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_245_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_66_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_122_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_61_seb);
  assign and_1735_nl = (nor_624_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[6]))
      & (fsm_output[1:0]==2'b11);
  assign mux_643_nl = MUX_s_1_2_2(and_1698_cse, and_1735_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm);
  assign nor_626_nl = ~((fsm_output[3:2]!=2'b00) | mux_643_nl);
  assign mux_644_nl = MUX_s_1_2_2(nor_626_nl, and_1669_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_260_nl = (mux_644_nl
      | or_dcpl_368) & and_220_ssc;
  assign and_1285_nl = (nor_624_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_14_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_itm))
      & and_dcpl_497 & and_220_ssc;
  assign mux_645_nl = MUX_s_1_2_2(nor_136_cse, and_1669_cse, fsm_output[4]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_62_nl
      = ~((~ MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_124_nl
      = MUX1HOT_v_5_3_2((MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_63_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_62_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_249_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_65_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_124_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_62_seb);
  assign and_1734_nl = (nor_620_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6]))
      & (fsm_output[1:0]==2'b11);
  assign mux_640_nl = MUX_s_1_2_2(and_1698_cse, and_1734_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm);
  assign nor_622_nl = ~((fsm_output[4:2]!=3'b000) | mux_640_nl);
  assign mux_641_nl = MUX_s_1_2_2(nor_622_nl, or_1113_cse, fsm_output[5]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_259_nl = (mux_641_nl
      | or_dcpl_150) & and_221_ssc;
  assign and_1281_nl = (nor_620_cse | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_16_tmp[6])
      | (~ ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_itm))
      & and_dcpl_497 & and_221_ssc;
  assign mux_642_nl = MUX_s_1_2_2(and_dcpl_223, or_1113_cse, fsm_output[5]);
  assign nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_1_sva_1[6:4])
      + 3'b001;
  assign MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[2:0];
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_34_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_34_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_35_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_35_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_36_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_36_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_37_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_37_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_38_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_38_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_39_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_39_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_40_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_40_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_41_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_41_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_42_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_42_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_43_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_43_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_44_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_44_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_45_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_45_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_46_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_46_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_47_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_47_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_48_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_48_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_49_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_49_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_50_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_50_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_51_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_51_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_52_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_52_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_53_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_53_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_54_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_54_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_55_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_55_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_56_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_56_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_57_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_57_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_58_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_58_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_59_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_59_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_60_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_60_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_61_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_61_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_62_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_62_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_63_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_63_sva_mx0w1[6:4])
      + 3'b001;
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva
      = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_sva_1[6:4])
      + 3'b001;
  assign MAC_3_r_ac_float_else_and_nl = MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_3_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_3_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_3_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva 
      = conv_s2s_6_7({MAC_3_r_ac_float_else_and_nl , MAC_3_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign mux_260_nl = MUX_s_1_2_2((fsm_output[1]), (~ or_dcpl_127), fsm_output[2]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_63_nl
      = ~((~ MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1)
      | (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2]));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_126_nl
      = MUX1HOT_v_5_3_2((MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_acc_sdt[4:0]),
      5'b10000, (MAC_64_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_acc_sdt[4:0]),
      {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_63_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_253_ssc , (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_psp_sva[2])});
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_64_nl
      = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux1h_126_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_63_seb);
  assign mux_261_nl = MUX_s_1_2_2(not_tmp_273, nor_tmp_66, fsm_output[7]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_nor_nl
      = ~(mux_261_nl | (fsm_output[8]));
  assign mux_559_nl = MUX_s_1_2_2(not_tmp_640, nor_tmp_66, fsm_output[7]);
  assign MAC_11_r_ac_float_else_and_nl = MUX_v_2_2_2(2'b00, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_1,
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign MAC_11_r_ac_float_else_and_1_nl = MUX_v_4_2_2(4'b0000, operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2,
      MAC_11_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_11_r_ac_float_else_and_nl , MAC_11_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_12_r_ac_float_else_and_nl = MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_12_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_12_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_12_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_12_r_ac_float_else_and_nl , MAC_12_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_13_r_ac_float_else_and_nl = MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_13_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_13_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_13_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_13_r_ac_float_else_and_nl , MAC_13_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_14_r_ac_float_else_and_nl = MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_14_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_14_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_14_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_14_r_ac_float_else_and_nl , MAC_14_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_15_r_ac_float_else_and_nl = MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_15_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_15_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_15_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_15_r_ac_float_else_and_nl , MAC_15_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_16_r_ac_float_else_and_nl = MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_16_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_16_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_16_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_16_r_ac_float_else_and_nl , MAC_16_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_17_r_ac_float_else_and_nl = MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_17_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_17_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_17_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_17_r_ac_float_else_and_nl , MAC_17_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_18_r_ac_float_else_and_nl = MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_18_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_18_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_18_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_18_r_ac_float_else_and_nl , MAC_18_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_19_r_ac_float_else_and_nl = MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_19_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_19_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_19_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_19_r_ac_float_else_and_nl , MAC_19_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_2_r_ac_float_else_and_nl = MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_2_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_2_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_2_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_2_r_ac_float_else_and_nl , MAC_2_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_20_r_ac_float_else_and_nl = MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_20_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_20_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_20_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_20_r_ac_float_else_and_nl , MAC_20_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_21_r_ac_float_else_and_nl = MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_21_r_ac_float_else_and_1_nl = MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      & MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_21_r_ac_float_else_and_2_nl = MUX_v_4_2_2(4'b0000, MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1,
      MAC_21_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_21_r_ac_float_else_and_nl , MAC_21_r_ac_float_else_and_1_nl
      , MAC_21_r_ac_float_else_and_2_nl}) + 7'b0000001;
  assign MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_22_r_ac_float_else_and_nl = MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_22_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_22_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_22_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_22_r_ac_float_else_and_nl , MAC_22_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_23_r_ac_float_else_and_nl = MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_23_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_23_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_23_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_23_r_ac_float_else_and_nl , MAC_23_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_24_r_ac_float_else_and_nl = MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_24_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_24_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_24_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_24_r_ac_float_else_and_nl , MAC_24_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_25_r_ac_float_else_and_nl = MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_25_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_25_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_25_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_25_r_ac_float_else_and_nl , MAC_25_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_26_r_ac_float_else_and_nl = MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_26_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_26_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_26_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_26_r_ac_float_else_and_nl , MAC_26_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_27_r_ac_float_else_and_nl = MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_27_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_27_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_27_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_27_r_ac_float_else_and_nl , MAC_27_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_28_r_ac_float_else_and_nl = MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_28_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_28_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_28_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_28_r_ac_float_else_and_nl , MAC_28_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_29_r_ac_float_else_and_nl = MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_29_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_29_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_29_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_29_r_ac_float_else_and_nl , MAC_29_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_30_r_ac_float_else_and_nl = MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_30_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_30_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_30_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_30_r_ac_float_else_and_nl , MAC_30_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_31_r_ac_float_else_and_nl = MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_31_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_31_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_31_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_31_r_ac_float_else_and_nl , MAC_31_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_32_r_ac_float_else_and_nl = MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_32_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_32_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_32_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_32_r_ac_float_else_and_nl , MAC_32_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_33_r_ac_float_else_and_nl = MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_5
      & MAC_33_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_33_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, MAC_33_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0,
      MAC_33_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_33_r_ac_float_else_and_nl , MAC_33_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_4_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_5
      & MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_4_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_43_lpi_1_dfm_4_0,
      MAC_4_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_4_r_ac_float_else_and_nl , MAC_4_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_5_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_5
      & MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_5_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_54_lpi_1_dfm_4_0,
      MAC_5_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_5_r_ac_float_else_and_nl , MAC_5_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_6_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_5
      & MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_6_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_60_lpi_1_dfm_4_0,
      MAC_6_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_6_r_ac_float_else_and_nl , MAC_6_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_7_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_5
      & MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_7_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_61_lpi_1_dfm_4_0,
      MAC_7_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_7_r_ac_float_else_and_nl , MAC_7_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_8_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_5
      & MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_8_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_62_lpi_1_dfm_4_0,
      MAC_8_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_8_r_ac_float_else_and_nl , MAC_8_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_9_r_ac_float_else_and_nl = ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_5
      & MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm;
  assign MAC_9_r_ac_float_else_and_1_nl = MUX_v_5_2_2(5'b00000, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_qr_6_0_63_lpi_1_dfm_4_0,
      MAC_9_r_ac_float_else_r_ac_float_else_r_ac_float_else_or_itm);
  assign nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl =
      conv_s2s_6_7({MAC_9_r_ac_float_else_and_nl , MAC_9_r_ac_float_else_and_1_nl})
      + 7'b0000001;
  assign MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl = nl_MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_nl[6:0];
  assign MAC_19_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_19_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_33_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_33_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_34_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_34_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_35_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_35_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_36_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_36_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_37_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_37_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_38_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_38_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_11_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_11_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_12_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_12_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_13_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_13_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_14_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_14_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_15_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_15_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_16_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_16_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_17_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_17_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_18_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_18_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_20_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_20_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_21_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_21_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_22_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_22_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_23_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_23_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_24_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_24_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_25_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_25_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_26_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_26_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_27_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_27_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_28_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_28_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_29_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_29_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_30_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_30_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_4_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_4_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_31_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_31_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign MAC_32_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_32_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_32_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_33_sva[21]))
      & MAC_33_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_59_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_59_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_31_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_32_sva[21]))
      & MAC_32_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_58_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_58_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_30_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_31_sva[21]))
      & MAC_31_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_57_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_57_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_29_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_30_sva[21]))
      & MAC_30_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_55_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_55_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_28_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_29_sva[21]))
      & MAC_29_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_54_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_54_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_27_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_28_sva[21]))
      & MAC_28_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_53_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_53_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_26_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_27_sva[21]))
      & MAC_27_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_52_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_52_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_25_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_26_sva[21]))
      & MAC_26_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_51_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_51_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_24_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_25_sva[21]))
      & MAC_25_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_6_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_6_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_23_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_24_sva[21]))
      & MAC_24_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_50_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_50_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_22_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_23_sva[21]))
      & MAC_23_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_49_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_49_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_21_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_22_sva[21]))
      & MAC_22_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_48_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_48_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_20_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_21_sva[21]))
      & MAC_21_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_47_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_47_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_19_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_20_sva[21]))
      & MAC_20_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_46_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_46_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_18_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_19_sva[21]))
      & MAC_19_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_45_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_45_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_17_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_18_sva[21]))
      & MAC_18_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_44_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_44_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_16_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_17_sva[21]))
      & MAC_17_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_43_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_43_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_15_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_16_sva[21]))
      & MAC_16_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_42_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_42_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_14_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_15_sva[21]))
      & MAC_15_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_41_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_41_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_13_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_14_sva[21]))
      & MAC_14_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_5_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_5_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_12_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_13_sva[21]))
      & MAC_13_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_11_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_12_sva[21]))
      & MAC_12_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_39_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_39_lpi_1_dfm_mx0w2!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_10_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_11_sva[21]))
      & MAC_11_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_2_nl
      = ~(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_all_sign_4_sva
      & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_3_sva[21])) & MAC_3_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_9_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_10_sva[21]))
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_12_itm);
  assign MAC_8_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_8_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_8_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_9_sva[21]))
      & MAC_9_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_63_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_63_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_7_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_8_sva[21]))
      & MAC_8_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_62_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_62_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_6_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_7_sva[21]))
      & MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_61_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_61_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_5_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_6_sva[21]))
      & MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_7_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_7_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_4_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_5_sva[21]))
      & MAC_5_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_60_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_60_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_3_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_4_sva[21]))
      & MAC_4_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign MAC_56_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_56_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign MAC_9_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_9_lpi_1_dfm_mx0w1!=11'b00000000000));
  assign MAC_3_ac_float_cctor_operator_ac_float_cctor_operator_nor_nl = ~((MAC_ac_float_cctor_m_3_lpi_1_dfm_mx0w4!=11'b00000000000));
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_if_nand_51_nl
      = ~(leading_sign_13_1_1_0_680f7e8f1e1ee1d0bfbb1629740d3a321b2d_55 & (~ (operator_13_2_true_AC_TRN_AC_WRAP_rshift_psp_10_sva_6_0_rsp_2[0])));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nand_1_nl
      = ~(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same_oreg & (~ (ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_r_m_2_sva[21]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_if_nor_itm);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_nand_nl
      = ~((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1[5:4]==2'b01));
  assign nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_7_lpi_1_dfm_6_0[3:0]);
  assign MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_or_1_nl = ((~((MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_109) | result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_mux_101_itm_mx0c7;
  assign and_270_nl = MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & and_dcpl_109;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_op_lshift_and_1_nl = (MAC_6_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_109;
  assign nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5:4])
      + 2'b01;
  assign MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_1_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = (z_out_1[5:4]) + 2'b01;
  assign MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl
      = nl_MAC_2_result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_nl[1:0];
  assign ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_mux1h_64_nl = MUX1HOT_s_1_3_2((MAC_10_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_sdt[5]),
      (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_acc_psp_1_sva_mx0w1[5]), (z_out_1[5]),
      {and_dcpl_105 , and_dcpl_154 , and_dcpl_157});
  assign nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl = nl_MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign nl_MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl
      = (~ (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]))
      + 5'b00001;
  assign MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl =
      nl_MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl[4:0];
  assign and_1310_nl = (~ (fsm_output[8])) & (fsm_output[2]) & (~ (fsm_output[3]))
      & and_dcpl_85 & and_dcpl_1276 & (~ (fsm_output[6])) & (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp
      | (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[5:4]!=2'b01));
  assign nand_55_nl = ~((fsm_output[1]) & or_351_cse);
  assign or_1170_nl = (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp
      & (fsm_output[2])) | (fsm_output[7:3]!=5'b00000);
  assign nor_645_nl = ~((~ result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_unequal_tmp)
      | (fsm_output[7:2]!=6'b000001));
  assign mux_658_nl = MUX_s_1_2_2(or_1170_nl, nor_645_nl, ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_11_sva);
  assign mux_659_nl = MUX_s_1_2_2(or_351_cse, mux_658_nl, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[4]);
  assign mux_660_nl = MUX_s_1_2_2(mux_659_nl, or_351_cse, result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_else_1_shift_l_mux_256_tmp[5]);
  assign or_1048_nl = (fsm_output[1]) | (~ mux_660_nl);
  assign mux_661_nl = MUX_s_1_2_2(nand_55_nl, or_1048_nl, fsm_output[0]);
  assign or_1565_nl = mux_661_nl | (fsm_output[8]);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_192_nl = (~ (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1312_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_193_nl = (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1312_m1c & (~ mux_1026_tmp);
  assign and_1315_nl = or_dcpl_308 & (~ (fsm_output[8])) & or_dcpl_105 & and_dcpl_1276;
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_194_nl = (~ (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1317_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_195_nl = (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1317_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_196_nl = (~ (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1318_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_197_nl = (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1318_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_198_nl = (~ (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1321_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_199_nl = (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1321_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_200_nl = (~ (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1322_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_201_nl = (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1322_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_202_nl = (~ (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1325_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_203_nl = (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1325_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_204_nl = (~ (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1326_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_205_nl = (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1326_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_206_nl = (~ (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1328_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_207_nl = (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1328_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_208_nl = (~ (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1329_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_209_nl = (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1329_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_210_nl = (~ (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1331_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_211_nl = (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1331_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_212_nl = (~ (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1332_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_213_nl = (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1332_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_214_nl = (~ (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1334_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_215_nl = (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1334_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_216_nl = (~ (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1335_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_217_nl = (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1335_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_218_nl = (~ (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1337_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_219_nl = (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1337_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_220_nl = (~ (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1338_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_221_nl = (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1338_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_222_nl = (~ (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1339_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_223_nl = (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1339_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_224_nl = (~ (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1340_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_225_nl = (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1340_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_226_nl = (~ (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1341_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_227_nl = (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1341_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_228_nl = (~ (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1342_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_229_nl = (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1342_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_230_nl = (~ (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1343_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_231_nl = (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1343_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_232_nl = (~ (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1344_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_233_nl = (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1344_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_234_nl = (~ (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1345_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_235_nl = (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1345_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_236_nl = (~ (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1346_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_237_nl = (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1346_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_238_nl = (~ (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1347_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_239_nl = (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1347_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_240_nl = (~ (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1348_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_241_nl = (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1348_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_242_nl = (~ (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1349_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_243_nl = (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1349_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_244_nl = (~ (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1350_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_245_nl = (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1350_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_246_nl = (~ (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1351_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_247_nl = (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1351_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_248_nl = (~ (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1352_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_249_nl = (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1352_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_250_nl = (~ (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1353_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_251_nl = (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1353_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_252_nl = (~ (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1354_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_253_nl = (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1354_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_254_nl = (~ (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1356_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_255_nl = (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1356_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_256_nl = (~ (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1357_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_257_nl = (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1357_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_258_nl = (~ (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1359_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_259_nl = (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1359_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_260_nl = (~ (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1360_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_261_nl = (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1360_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_262_nl = (~ (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1362_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_263_nl = (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1362_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_264_nl = (~ (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1363_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_265_nl = (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1363_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_266_nl = (~ (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1365_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_267_nl = (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1365_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_268_nl = (~ (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1366_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_269_nl = (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1366_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_270_nl = (~ (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1368_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_271_nl = (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1368_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_272_nl = (~ (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1369_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_273_nl = (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1369_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_274_nl = (~ (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1371_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_275_nl = (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1371_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_276_nl = (~ (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1372_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_277_nl = (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1372_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_278_nl = (~ (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1374_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_279_nl = (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1374_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_280_nl = (~ (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1375_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_281_nl = (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1375_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_282_nl = (~ (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1377_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_283_nl = (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1377_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_284_nl = (~ (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1378_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_285_nl = (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1378_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_286_nl = (~ (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1379_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_287_nl = (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1379_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_288_nl = (~ (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1380_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_289_nl = (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1380_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_290_nl = (~ (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1381_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_291_nl = (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1381_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_292_nl = (~ (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1382_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_293_nl = (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1382_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_294_nl = (~ (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1383_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_295_nl = (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1383_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_296_nl = (~ (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1384_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_297_nl = (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1384_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_298_nl = (~ (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1385_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_299_nl = (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1385_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_300_nl = (~ (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1386_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_301_nl = (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1386_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_302_nl = (~ (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1387_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_303_nl = (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1387_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_304_nl = (~ (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1388_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_305_nl = (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1388_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_306_nl = (~ (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1389_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_307_nl = (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1389_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_308_nl = (~ (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1390_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_309_nl = (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1390_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_310_nl = (~ (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1391_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_311_nl = (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1391_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_312_nl = (~ (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1392_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_313_nl = (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1392_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_314_nl = (~ (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1393_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_315_nl = (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1393_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_316_nl = (~ (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5]))
      & and_1394_m1c & (~ mux_1026_tmp);
  assign result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_317_nl = (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[5])
      & and_1394_m1c & (~ mux_1026_tmp);
  assign mux1h_1_nl = MUX1HOT_v_5_129_2((result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_1_lpi_1_dfm_1[4:0]),
      5'b01111, (MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_2_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_qr_5_0_3_lpi_1_dfm_1[4:0]),
      (MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_3_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_4_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_5_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_6_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_7_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_8_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]), MAC_9_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl,
      (MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_10_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_11_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_12_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_13_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_14_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_15_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_16_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_17_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_18_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_19_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_20_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_21_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_22_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_23_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_24_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_25_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_26_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_27_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_28_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_29_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_30_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_31_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_32_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_33_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_34_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_35_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_36_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_37_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_38_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_39_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_40_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_41_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_42_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_43_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_44_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_45_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_46_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_47_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_48_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_49_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_50_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_51_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_52_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_53_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_54_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_55_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_56_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_57_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_58_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_59_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_60_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_61_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_62_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_63_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, (MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_e_dif_acc_tmp[4:0]),
      MAC_64_result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_qelse_qif_acc_nl, {and_1310_nl
      , or_1565_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_192_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_193_nl
      , and_1315_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_194_nl ,
      result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_195_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_196_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_197_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_198_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_199_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_200_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_201_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_202_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_203_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_204_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_205_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_206_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_207_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_208_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_209_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_210_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_211_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_212_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_213_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_214_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_215_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_216_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_217_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_218_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_219_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_220_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_221_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_222_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_223_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_224_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_225_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_226_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_227_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_228_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_229_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_230_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_231_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_232_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_233_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_234_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_235_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_236_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_237_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_238_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_239_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_240_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_241_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_242_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_243_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_244_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_245_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_246_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_247_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_248_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_249_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_250_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_251_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_252_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_253_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_254_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_255_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_256_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_257_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_258_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_259_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_260_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_261_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_262_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_263_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_264_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_265_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_266_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_267_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_268_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_269_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_270_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_271_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_272_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_273_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_274_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_275_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_276_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_277_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_278_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_279_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_280_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_281_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_282_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_283_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_284_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_285_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_286_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_287_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_288_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_289_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_290_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_291_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_292_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_293_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_294_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_295_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_296_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_297_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_298_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_299_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_300_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_301_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_302_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_303_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_304_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_305_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_306_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_307_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_308_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_309_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_310_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_311_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_312_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_313_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_314_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_315_nl , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_316_nl
      , result_assign_from_n16_15_13_2_AC_TRN_AC_WRAP_and_317_nl});
  assign not_2129_nl = ~ mux_1026_tmp;
  assign and_1758_nl = MUX_v_5_2_2(5'b00000, mux1h_1_nl, not_2129_nl);
  assign nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      =  -(MAC_ac_float_cctor_m_8_lpi_1_dfm_6_0[3:0]);
  assign MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl
      = nl_MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_acc_nl[3:0];
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_nl = (~((MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      | MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1))
      & and_dcpl_109;
  assign and_272_nl = MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_shift_exponent_limited_acc_itm_6_1
      & (~ (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2]))
      & and_dcpl_109;
  assign result_plus_minus_11_1_5_AC_TRN_11_1_5_AC_TRN_add_r_and_1_nl = (MAC_7_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_actual_max_shift_left_acc_tmp[2])
      & and_dcpl_109;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl
      = MUX_v_7_2_2(MAC_ac_float_cctor_m_49_lpi_1_dfm_6_0, (signext_7_4(~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_acc_psp_3_sva[3:0]))),
      and_dcpl_1640);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl
      = ~(and_dcpl_1640 & (~(and_dcpl_1635 & (fsm_output[1:0]==2'b11) & and_dcpl_95)));
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_1_nl
      = ~(MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      | and_dcpl_1640);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      = MUX_v_4_2_2((~ MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1),
      4'b0001, and_dcpl_1640);
  assign nl_acc_nl = ({ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_3_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nand_1_nl})
      + conv_s2u_7_8({(~ and_dcpl_1640) , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_nor_1_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_else_1_qelse_mux_4_nl
      , 1'b1});
  assign acc_nl = nl_acc_nl[7:0];
  assign z_out = readslicef_8_7_1(acc_nl);
  assign and_1939_nl = or_351_cse & (~ (fsm_output[8])) & (fsm_output[0]) & (fsm_output[1]);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl
      = MUX_v_5_2_2((signext_5_4(~ (MAC_ac_float_cctor_m_62_lpi_1_dfm_6_0[3:0]))),
      ({MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_0
      , MAC_21_ac_float_11_1_5_AC_TRN_operator_11_1_5_AC_TRN_acc_1_itm_4_0_rsp_1}),
      and_1939_nl);
  assign nl_z_out_1 = conv_s2u_5_6(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_1_shift_r_mux_1_nl)
      + 6'b000001;
  assign z_out_1 = nl_z_out_1[5:0];
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_97_m1c = MUX_s_1_2_2((~
      MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1),
      (~ MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1),
      and_dcpl_1663);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_322_nl = (~ and_dcpl_1663)
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_97_m1c;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_323_nl = and_dcpl_1663
      & ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_97_m1c;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_318_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[10]))
      & MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_319_nl = (~ (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10]))
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_98_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_318_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_319_nl, and_dcpl_1663);
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_320_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva[10])
      & MAC_40_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_321_nl = (ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva[10])
      & MAC_2_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_if_3_nor_svs_1;
  assign ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_99_nl = MUX_s_1_2_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_320_nl,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_321_nl, and_dcpl_1663);
  assign z_out_2 = MUX1HOT_v_11_4_2(ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_40_sva,
      ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_op2_21_11_1_sva, 11'b01111111111,
      11'b10000000000, {ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_322_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_and_323_nl , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_98_nl
      , ac_float_cctor_assign_from_n32_31_22_2_AC_TRN_AC_WRAP_mux_99_nl});

  function automatic  MUX1HOT_s_1_129_2;
    input  input_128;
    input  input_127;
    input  input_126;
    input  input_125;
    input  input_124;
    input  input_123;
    input  input_122;
    input  input_121;
    input  input_120;
    input  input_119;
    input  input_118;
    input  input_117;
    input  input_116;
    input  input_115;
    input  input_114;
    input  input_113;
    input  input_112;
    input  input_111;
    input  input_110;
    input  input_109;
    input  input_108;
    input  input_107;
    input  input_106;
    input  input_105;
    input  input_104;
    input  input_103;
    input  input_102;
    input  input_101;
    input  input_100;
    input  input_99;
    input  input_98;
    input  input_97;
    input  input_96;
    input  input_95;
    input  input_94;
    input  input_93;
    input  input_92;
    input  input_91;
    input  input_90;
    input  input_89;
    input  input_88;
    input  input_87;
    input  input_86;
    input  input_85;
    input  input_84;
    input  input_83;
    input  input_82;
    input  input_81;
    input  input_80;
    input  input_79;
    input  input_78;
    input  input_77;
    input  input_76;
    input  input_75;
    input  input_74;
    input  input_73;
    input  input_72;
    input  input_71;
    input  input_70;
    input  input_69;
    input  input_68;
    input  input_67;
    input  input_66;
    input  input_65;
    input  input_64;
    input  input_63;
    input  input_62;
    input  input_61;
    input  input_60;
    input  input_59;
    input  input_58;
    input  input_57;
    input  input_56;
    input  input_55;
    input  input_54;
    input  input_53;
    input  input_52;
    input  input_51;
    input  input_50;
    input  input_49;
    input  input_48;
    input  input_47;
    input  input_46;
    input  input_45;
    input  input_44;
    input  input_43;
    input  input_42;
    input  input_41;
    input  input_40;
    input  input_39;
    input  input_38;
    input  input_37;
    input  input_36;
    input  input_35;
    input  input_34;
    input  input_33;
    input  input_32;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [128:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    result = result | (input_32 & sel[32]);
    result = result | (input_33 & sel[33]);
    result = result | (input_34 & sel[34]);
    result = result | (input_35 & sel[35]);
    result = result | (input_36 & sel[36]);
    result = result | (input_37 & sel[37]);
    result = result | (input_38 & sel[38]);
    result = result | (input_39 & sel[39]);
    result = result | (input_40 & sel[40]);
    result = result | (input_41 & sel[41]);
    result = result | (input_42 & sel[42]);
    result = result | (input_43 & sel[43]);
    result = result | (input_44 & sel[44]);
    result = result | (input_45 & sel[45]);
    result = result | (input_46 & sel[46]);
    result = result | (input_47 & sel[47]);
    result = result | (input_48 & sel[48]);
    result = result | (input_49 & sel[49]);
    result = result | (input_50 & sel[50]);
    result = result | (input_51 & sel[51]);
    result = result | (input_52 & sel[52]);
    result = result | (input_53 & sel[53]);
    result = result | (input_54 & sel[54]);
    result = result | (input_55 & sel[55]);
    result = result | (input_56 & sel[56]);
    result = result | (input_57 & sel[57]);
    result = result | (input_58 & sel[58]);
    result = result | (input_59 & sel[59]);
    result = result | (input_60 & sel[60]);
    result = result | (input_61 & sel[61]);
    result = result | (input_62 & sel[62]);
    result = result | (input_63 & sel[63]);
    result = result | (input_64 & sel[64]);
    result = result | (input_65 & sel[65]);
    result = result | (input_66 & sel[66]);
    result = result | (input_67 & sel[67]);
    result = result | (input_68 & sel[68]);
    result = result | (input_69 & sel[69]);
    result = result | (input_70 & sel[70]);
    result = result | (input_71 & sel[71]);
    result = result | (input_72 & sel[72]);
    result = result | (input_73 & sel[73]);
    result = result | (input_74 & sel[74]);
    result = result | (input_75 & sel[75]);
    result = result | (input_76 & sel[76]);
    result = result | (input_77 & sel[77]);
    result = result | (input_78 & sel[78]);
    result = result | (input_79 & sel[79]);
    result = result | (input_80 & sel[80]);
    result = result | (input_81 & sel[81]);
    result = result | (input_82 & sel[82]);
    result = result | (input_83 & sel[83]);
    result = result | (input_84 & sel[84]);
    result = result | (input_85 & sel[85]);
    result = result | (input_86 & sel[86]);
    result = result | (input_87 & sel[87]);
    result = result | (input_88 & sel[88]);
    result = result | (input_89 & sel[89]);
    result = result | (input_90 & sel[90]);
    result = result | (input_91 & sel[91]);
    result = result | (input_92 & sel[92]);
    result = result | (input_93 & sel[93]);
    result = result | (input_94 & sel[94]);
    result = result | (input_95 & sel[95]);
    result = result | (input_96 & sel[96]);
    result = result | (input_97 & sel[97]);
    result = result | (input_98 & sel[98]);
    result = result | (input_99 & sel[99]);
    result = result | (input_100 & sel[100]);
    result = result | (input_101 & sel[101]);
    result = result | (input_102 & sel[102]);
    result = result | (input_103 & sel[103]);
    result = result | (input_104 & sel[104]);
    result = result | (input_105 & sel[105]);
    result = result | (input_106 & sel[106]);
    result = result | (input_107 & sel[107]);
    result = result | (input_108 & sel[108]);
    result = result | (input_109 & sel[109]);
    result = result | (input_110 & sel[110]);
    result = result | (input_111 & sel[111]);
    result = result | (input_112 & sel[112]);
    result = result | (input_113 & sel[113]);
    result = result | (input_114 & sel[114]);
    result = result | (input_115 & sel[115]);
    result = result | (input_116 & sel[116]);
    result = result | (input_117 & sel[117]);
    result = result | (input_118 & sel[118]);
    result = result | (input_119 & sel[119]);
    result = result | (input_120 & sel[120]);
    result = result | (input_121 & sel[121]);
    result = result | (input_122 & sel[122]);
    result = result | (input_123 & sel[123]);
    result = result | (input_124 & sel[124]);
    result = result | (input_125 & sel[125]);
    result = result | (input_126 & sel[126]);
    result = result | (input_127 & sel[127]);
    result = result | (input_128 & sel[128]);
    MUX1HOT_s_1_129_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_3_2;
    input  input_2;
    input  input_1;
    input  input_0;
    input [2:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_4_2;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [3:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_5_2;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [4:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    MUX1HOT_s_1_5_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_64_2;
    input  input_63;
    input  input_62;
    input  input_61;
    input  input_60;
    input  input_59;
    input  input_58;
    input  input_57;
    input  input_56;
    input  input_55;
    input  input_54;
    input  input_53;
    input  input_52;
    input  input_51;
    input  input_50;
    input  input_49;
    input  input_48;
    input  input_47;
    input  input_46;
    input  input_45;
    input  input_44;
    input  input_43;
    input  input_42;
    input  input_41;
    input  input_40;
    input  input_39;
    input  input_38;
    input  input_37;
    input  input_36;
    input  input_35;
    input  input_34;
    input  input_33;
    input  input_32;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [63:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    result = result | (input_32 & sel[32]);
    result = result | (input_33 & sel[33]);
    result = result | (input_34 & sel[34]);
    result = result | (input_35 & sel[35]);
    result = result | (input_36 & sel[36]);
    result = result | (input_37 & sel[37]);
    result = result | (input_38 & sel[38]);
    result = result | (input_39 & sel[39]);
    result = result | (input_40 & sel[40]);
    result = result | (input_41 & sel[41]);
    result = result | (input_42 & sel[42]);
    result = result | (input_43 & sel[43]);
    result = result | (input_44 & sel[44]);
    result = result | (input_45 & sel[45]);
    result = result | (input_46 & sel[46]);
    result = result | (input_47 & sel[47]);
    result = result | (input_48 & sel[48]);
    result = result | (input_49 & sel[49]);
    result = result | (input_50 & sel[50]);
    result = result | (input_51 & sel[51]);
    result = result | (input_52 & sel[52]);
    result = result | (input_53 & sel[53]);
    result = result | (input_54 & sel[54]);
    result = result | (input_55 & sel[55]);
    result = result | (input_56 & sel[56]);
    result = result | (input_57 & sel[57]);
    result = result | (input_58 & sel[58]);
    result = result | (input_59 & sel[59]);
    result = result | (input_60 & sel[60]);
    result = result | (input_61 & sel[61]);
    result = result | (input_62 & sel[62]);
    result = result | (input_63 & sel[63]);
    MUX1HOT_s_1_64_2 = result;
  end
  endfunction


  function automatic  MUX1HOT_s_1_67_2;
    input  input_66;
    input  input_65;
    input  input_64;
    input  input_63;
    input  input_62;
    input  input_61;
    input  input_60;
    input  input_59;
    input  input_58;
    input  input_57;
    input  input_56;
    input  input_55;
    input  input_54;
    input  input_53;
    input  input_52;
    input  input_51;
    input  input_50;
    input  input_49;
    input  input_48;
    input  input_47;
    input  input_46;
    input  input_45;
    input  input_44;
    input  input_43;
    input  input_42;
    input  input_41;
    input  input_40;
    input  input_39;
    input  input_38;
    input  input_37;
    input  input_36;
    input  input_35;
    input  input_34;
    input  input_33;
    input  input_32;
    input  input_31;
    input  input_30;
    input  input_29;
    input  input_28;
    input  input_27;
    input  input_26;
    input  input_25;
    input  input_24;
    input  input_23;
    input  input_22;
    input  input_21;
    input  input_20;
    input  input_19;
    input  input_18;
    input  input_17;
    input  input_16;
    input  input_15;
    input  input_14;
    input  input_13;
    input  input_12;
    input  input_11;
    input  input_10;
    input  input_9;
    input  input_8;
    input  input_7;
    input  input_6;
    input  input_5;
    input  input_4;
    input  input_3;
    input  input_2;
    input  input_1;
    input  input_0;
    input [66:0] sel;
    reg  result;
  begin
    result = input_0 & sel[0];
    result = result | (input_1 & sel[1]);
    result = result | (input_2 & sel[2]);
    result = result | (input_3 & sel[3]);
    result = result | (input_4 & sel[4]);
    result = result | (input_5 & sel[5]);
    result = result | (input_6 & sel[6]);
    result = result | (input_7 & sel[7]);
    result = result | (input_8 & sel[8]);
    result = result | (input_9 & sel[9]);
    result = result | (input_10 & sel[10]);
    result = result | (input_11 & sel[11]);
    result = result | (input_12 & sel[12]);
    result = result | (input_13 & sel[13]);
    result = result | (input_14 & sel[14]);
    result = result | (input_15 & sel[15]);
    result = result | (input_16 & sel[16]);
    result = result | (input_17 & sel[17]);
    result = result | (input_18 & sel[18]);
    result = result | (input_19 & sel[19]);
    result = result | (input_20 & sel[20]);
    result = result | (input_21 & sel[21]);
    result = result | (input_22 & sel[22]);
    result = result | (input_23 & sel[23]);
    result = result | (input_24 & sel[24]);
    result = result | (input_25 & sel[25]);
    result = result | (input_26 & sel[26]);
    result = result | (input_27 & sel[27]);
    result = result | (input_28 & sel[28]);
    result = result | (input_29 & sel[29]);
    result = result | (input_30 & sel[30]);
    result = result | (input_31 & sel[31]);
    result = result | (input_32 & sel[32]);
    result = result | (input_33 & sel[33]);
    result = result | (input_34 & sel[34]);
    result = result | (input_35 & sel[35]);
    result = result | (input_36 & sel[36]);
    result = result | (input_37 & sel[37]);
    result = result | (input_38 & sel[38]);
    result = result | (input_39 & sel[39]);
    result = result | (input_40 & sel[40]);
    result = result | (input_41 & sel[41]);
    result = result | (input_42 & sel[42]);
    result = result | (input_43 & sel[43]);
    result = result | (input_44 & sel[44]);
    result = result | (input_45 & sel[45]);
    result = result | (input_46 & sel[46]);
    result = result | (input_47 & sel[47]);
    result = result | (input_48 & sel[48]);
    result = result | (input_49 & sel[49]);
    result = result | (input_50 & sel[50]);
    result = result | (input_51 & sel[51]);
    result = result | (input_52 & sel[52]);
    result = result | (input_53 & sel[53]);
    result = result | (input_54 & sel[54]);
    result = result | (input_55 & sel[55]);
    result = result | (input_56 & sel[56]);
    result = result | (input_57 & sel[57]);
    result = result | (input_58 & sel[58]);
    result = result | (input_59 & sel[59]);
    result = result | (input_60 & sel[60]);
    result = result | (input_61 & sel[61]);
    result = result | (input_62 & sel[62]);
    result = result | (input_63 & sel[63]);
    result = result | (input_64 & sel[64]);
    result = result | (input_65 & sel[65]);
    result = result | (input_66 & sel[66]);
    MUX1HOT_s_1_67_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_3_2;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [2:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    MUX1HOT_v_11_3_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_4_2;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [3:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    MUX1HOT_v_11_4_2 = result;
  end
  endfunction


  function automatic [10:0] MUX1HOT_v_11_5_2;
    input [10:0] input_4;
    input [10:0] input_3;
    input [10:0] input_2;
    input [10:0] input_1;
    input [10:0] input_0;
    input [4:0] sel;
    reg [10:0] result;
  begin
    result = input_0 & {11{sel[0]}};
    result = result | (input_1 & {11{sel[1]}});
    result = result | (input_2 & {11{sel[2]}});
    result = result | (input_3 & {11{sel[3]}});
    result = result | (input_4 & {11{sel[4]}});
    MUX1HOT_v_11_5_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_130_2;
    input [1:0] input_129;
    input [1:0] input_128;
    input [1:0] input_127;
    input [1:0] input_126;
    input [1:0] input_125;
    input [1:0] input_124;
    input [1:0] input_123;
    input [1:0] input_122;
    input [1:0] input_121;
    input [1:0] input_120;
    input [1:0] input_119;
    input [1:0] input_118;
    input [1:0] input_117;
    input [1:0] input_116;
    input [1:0] input_115;
    input [1:0] input_114;
    input [1:0] input_113;
    input [1:0] input_112;
    input [1:0] input_111;
    input [1:0] input_110;
    input [1:0] input_109;
    input [1:0] input_108;
    input [1:0] input_107;
    input [1:0] input_106;
    input [1:0] input_105;
    input [1:0] input_104;
    input [1:0] input_103;
    input [1:0] input_102;
    input [1:0] input_101;
    input [1:0] input_100;
    input [1:0] input_99;
    input [1:0] input_98;
    input [1:0] input_97;
    input [1:0] input_96;
    input [1:0] input_95;
    input [1:0] input_94;
    input [1:0] input_93;
    input [1:0] input_92;
    input [1:0] input_91;
    input [1:0] input_90;
    input [1:0] input_89;
    input [1:0] input_88;
    input [1:0] input_87;
    input [1:0] input_86;
    input [1:0] input_85;
    input [1:0] input_84;
    input [1:0] input_83;
    input [1:0] input_82;
    input [1:0] input_81;
    input [1:0] input_80;
    input [1:0] input_79;
    input [1:0] input_78;
    input [1:0] input_77;
    input [1:0] input_76;
    input [1:0] input_75;
    input [1:0] input_74;
    input [1:0] input_73;
    input [1:0] input_72;
    input [1:0] input_71;
    input [1:0] input_70;
    input [1:0] input_69;
    input [1:0] input_68;
    input [1:0] input_67;
    input [1:0] input_66;
    input [1:0] input_65;
    input [1:0] input_64;
    input [1:0] input_63;
    input [1:0] input_62;
    input [1:0] input_61;
    input [1:0] input_60;
    input [1:0] input_59;
    input [1:0] input_58;
    input [1:0] input_57;
    input [1:0] input_56;
    input [1:0] input_55;
    input [1:0] input_54;
    input [1:0] input_53;
    input [1:0] input_52;
    input [1:0] input_51;
    input [1:0] input_50;
    input [1:0] input_49;
    input [1:0] input_48;
    input [1:0] input_47;
    input [1:0] input_46;
    input [1:0] input_45;
    input [1:0] input_44;
    input [1:0] input_43;
    input [1:0] input_42;
    input [1:0] input_41;
    input [1:0] input_40;
    input [1:0] input_39;
    input [1:0] input_38;
    input [1:0] input_37;
    input [1:0] input_36;
    input [1:0] input_35;
    input [1:0] input_34;
    input [1:0] input_33;
    input [1:0] input_32;
    input [1:0] input_31;
    input [1:0] input_30;
    input [1:0] input_29;
    input [1:0] input_28;
    input [1:0] input_27;
    input [1:0] input_26;
    input [1:0] input_25;
    input [1:0] input_24;
    input [1:0] input_23;
    input [1:0] input_22;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [129:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    result = result | (input_22 & {2{sel[22]}});
    result = result | (input_23 & {2{sel[23]}});
    result = result | (input_24 & {2{sel[24]}});
    result = result | (input_25 & {2{sel[25]}});
    result = result | (input_26 & {2{sel[26]}});
    result = result | (input_27 & {2{sel[27]}});
    result = result | (input_28 & {2{sel[28]}});
    result = result | (input_29 & {2{sel[29]}});
    result = result | (input_30 & {2{sel[30]}});
    result = result | (input_31 & {2{sel[31]}});
    result = result | (input_32 & {2{sel[32]}});
    result = result | (input_33 & {2{sel[33]}});
    result = result | (input_34 & {2{sel[34]}});
    result = result | (input_35 & {2{sel[35]}});
    result = result | (input_36 & {2{sel[36]}});
    result = result | (input_37 & {2{sel[37]}});
    result = result | (input_38 & {2{sel[38]}});
    result = result | (input_39 & {2{sel[39]}});
    result = result | (input_40 & {2{sel[40]}});
    result = result | (input_41 & {2{sel[41]}});
    result = result | (input_42 & {2{sel[42]}});
    result = result | (input_43 & {2{sel[43]}});
    result = result | (input_44 & {2{sel[44]}});
    result = result | (input_45 & {2{sel[45]}});
    result = result | (input_46 & {2{sel[46]}});
    result = result | (input_47 & {2{sel[47]}});
    result = result | (input_48 & {2{sel[48]}});
    result = result | (input_49 & {2{sel[49]}});
    result = result | (input_50 & {2{sel[50]}});
    result = result | (input_51 & {2{sel[51]}});
    result = result | (input_52 & {2{sel[52]}});
    result = result | (input_53 & {2{sel[53]}});
    result = result | (input_54 & {2{sel[54]}});
    result = result | (input_55 & {2{sel[55]}});
    result = result | (input_56 & {2{sel[56]}});
    result = result | (input_57 & {2{sel[57]}});
    result = result | (input_58 & {2{sel[58]}});
    result = result | (input_59 & {2{sel[59]}});
    result = result | (input_60 & {2{sel[60]}});
    result = result | (input_61 & {2{sel[61]}});
    result = result | (input_62 & {2{sel[62]}});
    result = result | (input_63 & {2{sel[63]}});
    result = result | (input_64 & {2{sel[64]}});
    result = result | (input_65 & {2{sel[65]}});
    result = result | (input_66 & {2{sel[66]}});
    result = result | (input_67 & {2{sel[67]}});
    result = result | (input_68 & {2{sel[68]}});
    result = result | (input_69 & {2{sel[69]}});
    result = result | (input_70 & {2{sel[70]}});
    result = result | (input_71 & {2{sel[71]}});
    result = result | (input_72 & {2{sel[72]}});
    result = result | (input_73 & {2{sel[73]}});
    result = result | (input_74 & {2{sel[74]}});
    result = result | (input_75 & {2{sel[75]}});
    result = result | (input_76 & {2{sel[76]}});
    result = result | (input_77 & {2{sel[77]}});
    result = result | (input_78 & {2{sel[78]}});
    result = result | (input_79 & {2{sel[79]}});
    result = result | (input_80 & {2{sel[80]}});
    result = result | (input_81 & {2{sel[81]}});
    result = result | (input_82 & {2{sel[82]}});
    result = result | (input_83 & {2{sel[83]}});
    result = result | (input_84 & {2{sel[84]}});
    result = result | (input_85 & {2{sel[85]}});
    result = result | (input_86 & {2{sel[86]}});
    result = result | (input_87 & {2{sel[87]}});
    result = result | (input_88 & {2{sel[88]}});
    result = result | (input_89 & {2{sel[89]}});
    result = result | (input_90 & {2{sel[90]}});
    result = result | (input_91 & {2{sel[91]}});
    result = result | (input_92 & {2{sel[92]}});
    result = result | (input_93 & {2{sel[93]}});
    result = result | (input_94 & {2{sel[94]}});
    result = result | (input_95 & {2{sel[95]}});
    result = result | (input_96 & {2{sel[96]}});
    result = result | (input_97 & {2{sel[97]}});
    result = result | (input_98 & {2{sel[98]}});
    result = result | (input_99 & {2{sel[99]}});
    result = result | (input_100 & {2{sel[100]}});
    result = result | (input_101 & {2{sel[101]}});
    result = result | (input_102 & {2{sel[102]}});
    result = result | (input_103 & {2{sel[103]}});
    result = result | (input_104 & {2{sel[104]}});
    result = result | (input_105 & {2{sel[105]}});
    result = result | (input_106 & {2{sel[106]}});
    result = result | (input_107 & {2{sel[107]}});
    result = result | (input_108 & {2{sel[108]}});
    result = result | (input_109 & {2{sel[109]}});
    result = result | (input_110 & {2{sel[110]}});
    result = result | (input_111 & {2{sel[111]}});
    result = result | (input_112 & {2{sel[112]}});
    result = result | (input_113 & {2{sel[113]}});
    result = result | (input_114 & {2{sel[114]}});
    result = result | (input_115 & {2{sel[115]}});
    result = result | (input_116 & {2{sel[116]}});
    result = result | (input_117 & {2{sel[117]}});
    result = result | (input_118 & {2{sel[118]}});
    result = result | (input_119 & {2{sel[119]}});
    result = result | (input_120 & {2{sel[120]}});
    result = result | (input_121 & {2{sel[121]}});
    result = result | (input_122 & {2{sel[122]}});
    result = result | (input_123 & {2{sel[123]}});
    result = result | (input_124 & {2{sel[124]}});
    result = result | (input_125 & {2{sel[125]}});
    result = result | (input_126 & {2{sel[126]}});
    result = result | (input_127 & {2{sel[127]}});
    result = result | (input_128 & {2{sel[128]}});
    result = result | (input_129 & {2{sel[129]}});
    MUX1HOT_v_2_130_2 = result;
  end
  endfunction


  function automatic [1:0] MUX1HOT_v_2_64_2;
    input [1:0] input_63;
    input [1:0] input_62;
    input [1:0] input_61;
    input [1:0] input_60;
    input [1:0] input_59;
    input [1:0] input_58;
    input [1:0] input_57;
    input [1:0] input_56;
    input [1:0] input_55;
    input [1:0] input_54;
    input [1:0] input_53;
    input [1:0] input_52;
    input [1:0] input_51;
    input [1:0] input_50;
    input [1:0] input_49;
    input [1:0] input_48;
    input [1:0] input_47;
    input [1:0] input_46;
    input [1:0] input_45;
    input [1:0] input_44;
    input [1:0] input_43;
    input [1:0] input_42;
    input [1:0] input_41;
    input [1:0] input_40;
    input [1:0] input_39;
    input [1:0] input_38;
    input [1:0] input_37;
    input [1:0] input_36;
    input [1:0] input_35;
    input [1:0] input_34;
    input [1:0] input_33;
    input [1:0] input_32;
    input [1:0] input_31;
    input [1:0] input_30;
    input [1:0] input_29;
    input [1:0] input_28;
    input [1:0] input_27;
    input [1:0] input_26;
    input [1:0] input_25;
    input [1:0] input_24;
    input [1:0] input_23;
    input [1:0] input_22;
    input [1:0] input_21;
    input [1:0] input_20;
    input [1:0] input_19;
    input [1:0] input_18;
    input [1:0] input_17;
    input [1:0] input_16;
    input [1:0] input_15;
    input [1:0] input_14;
    input [1:0] input_13;
    input [1:0] input_12;
    input [1:0] input_11;
    input [1:0] input_10;
    input [1:0] input_9;
    input [1:0] input_8;
    input [1:0] input_7;
    input [1:0] input_6;
    input [1:0] input_5;
    input [1:0] input_4;
    input [1:0] input_3;
    input [1:0] input_2;
    input [1:0] input_1;
    input [1:0] input_0;
    input [63:0] sel;
    reg [1:0] result;
  begin
    result = input_0 & {2{sel[0]}};
    result = result | (input_1 & {2{sel[1]}});
    result = result | (input_2 & {2{sel[2]}});
    result = result | (input_3 & {2{sel[3]}});
    result = result | (input_4 & {2{sel[4]}});
    result = result | (input_5 & {2{sel[5]}});
    result = result | (input_6 & {2{sel[6]}});
    result = result | (input_7 & {2{sel[7]}});
    result = result | (input_8 & {2{sel[8]}});
    result = result | (input_9 & {2{sel[9]}});
    result = result | (input_10 & {2{sel[10]}});
    result = result | (input_11 & {2{sel[11]}});
    result = result | (input_12 & {2{sel[12]}});
    result = result | (input_13 & {2{sel[13]}});
    result = result | (input_14 & {2{sel[14]}});
    result = result | (input_15 & {2{sel[15]}});
    result = result | (input_16 & {2{sel[16]}});
    result = result | (input_17 & {2{sel[17]}});
    result = result | (input_18 & {2{sel[18]}});
    result = result | (input_19 & {2{sel[19]}});
    result = result | (input_20 & {2{sel[20]}});
    result = result | (input_21 & {2{sel[21]}});
    result = result | (input_22 & {2{sel[22]}});
    result = result | (input_23 & {2{sel[23]}});
    result = result | (input_24 & {2{sel[24]}});
    result = result | (input_25 & {2{sel[25]}});
    result = result | (input_26 & {2{sel[26]}});
    result = result | (input_27 & {2{sel[27]}});
    result = result | (input_28 & {2{sel[28]}});
    result = result | (input_29 & {2{sel[29]}});
    result = result | (input_30 & {2{sel[30]}});
    result = result | (input_31 & {2{sel[31]}});
    result = result | (input_32 & {2{sel[32]}});
    result = result | (input_33 & {2{sel[33]}});
    result = result | (input_34 & {2{sel[34]}});
    result = result | (input_35 & {2{sel[35]}});
    result = result | (input_36 & {2{sel[36]}});
    result = result | (input_37 & {2{sel[37]}});
    result = result | (input_38 & {2{sel[38]}});
    result = result | (input_39 & {2{sel[39]}});
    result = result | (input_40 & {2{sel[40]}});
    result = result | (input_41 & {2{sel[41]}});
    result = result | (input_42 & {2{sel[42]}});
    result = result | (input_43 & {2{sel[43]}});
    result = result | (input_44 & {2{sel[44]}});
    result = result | (input_45 & {2{sel[45]}});
    result = result | (input_46 & {2{sel[46]}});
    result = result | (input_47 & {2{sel[47]}});
    result = result | (input_48 & {2{sel[48]}});
    result = result | (input_49 & {2{sel[49]}});
    result = result | (input_50 & {2{sel[50]}});
    result = result | (input_51 & {2{sel[51]}});
    result = result | (input_52 & {2{sel[52]}});
    result = result | (input_53 & {2{sel[53]}});
    result = result | (input_54 & {2{sel[54]}});
    result = result | (input_55 & {2{sel[55]}});
    result = result | (input_56 & {2{sel[56]}});
    result = result | (input_57 & {2{sel[57]}});
    result = result | (input_58 & {2{sel[58]}});
    result = result | (input_59 & {2{sel[59]}});
    result = result | (input_60 & {2{sel[60]}});
    result = result | (input_61 & {2{sel[61]}});
    result = result | (input_62 & {2{sel[62]}});
    result = result | (input_63 & {2{sel[63]}});
    MUX1HOT_v_2_64_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_128_2;
    input [3:0] input_127;
    input [3:0] input_126;
    input [3:0] input_125;
    input [3:0] input_124;
    input [3:0] input_123;
    input [3:0] input_122;
    input [3:0] input_121;
    input [3:0] input_120;
    input [3:0] input_119;
    input [3:0] input_118;
    input [3:0] input_117;
    input [3:0] input_116;
    input [3:0] input_115;
    input [3:0] input_114;
    input [3:0] input_113;
    input [3:0] input_112;
    input [3:0] input_111;
    input [3:0] input_110;
    input [3:0] input_109;
    input [3:0] input_108;
    input [3:0] input_107;
    input [3:0] input_106;
    input [3:0] input_105;
    input [3:0] input_104;
    input [3:0] input_103;
    input [3:0] input_102;
    input [3:0] input_101;
    input [3:0] input_100;
    input [3:0] input_99;
    input [3:0] input_98;
    input [3:0] input_97;
    input [3:0] input_96;
    input [3:0] input_95;
    input [3:0] input_94;
    input [3:0] input_93;
    input [3:0] input_92;
    input [3:0] input_91;
    input [3:0] input_90;
    input [3:0] input_89;
    input [3:0] input_88;
    input [3:0] input_87;
    input [3:0] input_86;
    input [3:0] input_85;
    input [3:0] input_84;
    input [3:0] input_83;
    input [3:0] input_82;
    input [3:0] input_81;
    input [3:0] input_80;
    input [3:0] input_79;
    input [3:0] input_78;
    input [3:0] input_77;
    input [3:0] input_76;
    input [3:0] input_75;
    input [3:0] input_74;
    input [3:0] input_73;
    input [3:0] input_72;
    input [3:0] input_71;
    input [3:0] input_70;
    input [3:0] input_69;
    input [3:0] input_68;
    input [3:0] input_67;
    input [3:0] input_66;
    input [3:0] input_65;
    input [3:0] input_64;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [127:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    result = result | (input_51 & {4{sel[51]}});
    result = result | (input_52 & {4{sel[52]}});
    result = result | (input_53 & {4{sel[53]}});
    result = result | (input_54 & {4{sel[54]}});
    result = result | (input_55 & {4{sel[55]}});
    result = result | (input_56 & {4{sel[56]}});
    result = result | (input_57 & {4{sel[57]}});
    result = result | (input_58 & {4{sel[58]}});
    result = result | (input_59 & {4{sel[59]}});
    result = result | (input_60 & {4{sel[60]}});
    result = result | (input_61 & {4{sel[61]}});
    result = result | (input_62 & {4{sel[62]}});
    result = result | (input_63 & {4{sel[63]}});
    result = result | (input_64 & {4{sel[64]}});
    result = result | (input_65 & {4{sel[65]}});
    result = result | (input_66 & {4{sel[66]}});
    result = result | (input_67 & {4{sel[67]}});
    result = result | (input_68 & {4{sel[68]}});
    result = result | (input_69 & {4{sel[69]}});
    result = result | (input_70 & {4{sel[70]}});
    result = result | (input_71 & {4{sel[71]}});
    result = result | (input_72 & {4{sel[72]}});
    result = result | (input_73 & {4{sel[73]}});
    result = result | (input_74 & {4{sel[74]}});
    result = result | (input_75 & {4{sel[75]}});
    result = result | (input_76 & {4{sel[76]}});
    result = result | (input_77 & {4{sel[77]}});
    result = result | (input_78 & {4{sel[78]}});
    result = result | (input_79 & {4{sel[79]}});
    result = result | (input_80 & {4{sel[80]}});
    result = result | (input_81 & {4{sel[81]}});
    result = result | (input_82 & {4{sel[82]}});
    result = result | (input_83 & {4{sel[83]}});
    result = result | (input_84 & {4{sel[84]}});
    result = result | (input_85 & {4{sel[85]}});
    result = result | (input_86 & {4{sel[86]}});
    result = result | (input_87 & {4{sel[87]}});
    result = result | (input_88 & {4{sel[88]}});
    result = result | (input_89 & {4{sel[89]}});
    result = result | (input_90 & {4{sel[90]}});
    result = result | (input_91 & {4{sel[91]}});
    result = result | (input_92 & {4{sel[92]}});
    result = result | (input_93 & {4{sel[93]}});
    result = result | (input_94 & {4{sel[94]}});
    result = result | (input_95 & {4{sel[95]}});
    result = result | (input_96 & {4{sel[96]}});
    result = result | (input_97 & {4{sel[97]}});
    result = result | (input_98 & {4{sel[98]}});
    result = result | (input_99 & {4{sel[99]}});
    result = result | (input_100 & {4{sel[100]}});
    result = result | (input_101 & {4{sel[101]}});
    result = result | (input_102 & {4{sel[102]}});
    result = result | (input_103 & {4{sel[103]}});
    result = result | (input_104 & {4{sel[104]}});
    result = result | (input_105 & {4{sel[105]}});
    result = result | (input_106 & {4{sel[106]}});
    result = result | (input_107 & {4{sel[107]}});
    result = result | (input_108 & {4{sel[108]}});
    result = result | (input_109 & {4{sel[109]}});
    result = result | (input_110 & {4{sel[110]}});
    result = result | (input_111 & {4{sel[111]}});
    result = result | (input_112 & {4{sel[112]}});
    result = result | (input_113 & {4{sel[113]}});
    result = result | (input_114 & {4{sel[114]}});
    result = result | (input_115 & {4{sel[115]}});
    result = result | (input_116 & {4{sel[116]}});
    result = result | (input_117 & {4{sel[117]}});
    result = result | (input_118 & {4{sel[118]}});
    result = result | (input_119 & {4{sel[119]}});
    result = result | (input_120 & {4{sel[120]}});
    result = result | (input_121 & {4{sel[121]}});
    result = result | (input_122 & {4{sel[122]}});
    result = result | (input_123 & {4{sel[123]}});
    result = result | (input_124 & {4{sel[124]}});
    result = result | (input_125 & {4{sel[125]}});
    result = result | (input_126 & {4{sel[126]}});
    result = result | (input_127 & {4{sel[127]}});
    MUX1HOT_v_4_128_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_130_2;
    input [3:0] input_129;
    input [3:0] input_128;
    input [3:0] input_127;
    input [3:0] input_126;
    input [3:0] input_125;
    input [3:0] input_124;
    input [3:0] input_123;
    input [3:0] input_122;
    input [3:0] input_121;
    input [3:0] input_120;
    input [3:0] input_119;
    input [3:0] input_118;
    input [3:0] input_117;
    input [3:0] input_116;
    input [3:0] input_115;
    input [3:0] input_114;
    input [3:0] input_113;
    input [3:0] input_112;
    input [3:0] input_111;
    input [3:0] input_110;
    input [3:0] input_109;
    input [3:0] input_108;
    input [3:0] input_107;
    input [3:0] input_106;
    input [3:0] input_105;
    input [3:0] input_104;
    input [3:0] input_103;
    input [3:0] input_102;
    input [3:0] input_101;
    input [3:0] input_100;
    input [3:0] input_99;
    input [3:0] input_98;
    input [3:0] input_97;
    input [3:0] input_96;
    input [3:0] input_95;
    input [3:0] input_94;
    input [3:0] input_93;
    input [3:0] input_92;
    input [3:0] input_91;
    input [3:0] input_90;
    input [3:0] input_89;
    input [3:0] input_88;
    input [3:0] input_87;
    input [3:0] input_86;
    input [3:0] input_85;
    input [3:0] input_84;
    input [3:0] input_83;
    input [3:0] input_82;
    input [3:0] input_81;
    input [3:0] input_80;
    input [3:0] input_79;
    input [3:0] input_78;
    input [3:0] input_77;
    input [3:0] input_76;
    input [3:0] input_75;
    input [3:0] input_74;
    input [3:0] input_73;
    input [3:0] input_72;
    input [3:0] input_71;
    input [3:0] input_70;
    input [3:0] input_69;
    input [3:0] input_68;
    input [3:0] input_67;
    input [3:0] input_66;
    input [3:0] input_65;
    input [3:0] input_64;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [129:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    result = result | (input_51 & {4{sel[51]}});
    result = result | (input_52 & {4{sel[52]}});
    result = result | (input_53 & {4{sel[53]}});
    result = result | (input_54 & {4{sel[54]}});
    result = result | (input_55 & {4{sel[55]}});
    result = result | (input_56 & {4{sel[56]}});
    result = result | (input_57 & {4{sel[57]}});
    result = result | (input_58 & {4{sel[58]}});
    result = result | (input_59 & {4{sel[59]}});
    result = result | (input_60 & {4{sel[60]}});
    result = result | (input_61 & {4{sel[61]}});
    result = result | (input_62 & {4{sel[62]}});
    result = result | (input_63 & {4{sel[63]}});
    result = result | (input_64 & {4{sel[64]}});
    result = result | (input_65 & {4{sel[65]}});
    result = result | (input_66 & {4{sel[66]}});
    result = result | (input_67 & {4{sel[67]}});
    result = result | (input_68 & {4{sel[68]}});
    result = result | (input_69 & {4{sel[69]}});
    result = result | (input_70 & {4{sel[70]}});
    result = result | (input_71 & {4{sel[71]}});
    result = result | (input_72 & {4{sel[72]}});
    result = result | (input_73 & {4{sel[73]}});
    result = result | (input_74 & {4{sel[74]}});
    result = result | (input_75 & {4{sel[75]}});
    result = result | (input_76 & {4{sel[76]}});
    result = result | (input_77 & {4{sel[77]}});
    result = result | (input_78 & {4{sel[78]}});
    result = result | (input_79 & {4{sel[79]}});
    result = result | (input_80 & {4{sel[80]}});
    result = result | (input_81 & {4{sel[81]}});
    result = result | (input_82 & {4{sel[82]}});
    result = result | (input_83 & {4{sel[83]}});
    result = result | (input_84 & {4{sel[84]}});
    result = result | (input_85 & {4{sel[85]}});
    result = result | (input_86 & {4{sel[86]}});
    result = result | (input_87 & {4{sel[87]}});
    result = result | (input_88 & {4{sel[88]}});
    result = result | (input_89 & {4{sel[89]}});
    result = result | (input_90 & {4{sel[90]}});
    result = result | (input_91 & {4{sel[91]}});
    result = result | (input_92 & {4{sel[92]}});
    result = result | (input_93 & {4{sel[93]}});
    result = result | (input_94 & {4{sel[94]}});
    result = result | (input_95 & {4{sel[95]}});
    result = result | (input_96 & {4{sel[96]}});
    result = result | (input_97 & {4{sel[97]}});
    result = result | (input_98 & {4{sel[98]}});
    result = result | (input_99 & {4{sel[99]}});
    result = result | (input_100 & {4{sel[100]}});
    result = result | (input_101 & {4{sel[101]}});
    result = result | (input_102 & {4{sel[102]}});
    result = result | (input_103 & {4{sel[103]}});
    result = result | (input_104 & {4{sel[104]}});
    result = result | (input_105 & {4{sel[105]}});
    result = result | (input_106 & {4{sel[106]}});
    result = result | (input_107 & {4{sel[107]}});
    result = result | (input_108 & {4{sel[108]}});
    result = result | (input_109 & {4{sel[109]}});
    result = result | (input_110 & {4{sel[110]}});
    result = result | (input_111 & {4{sel[111]}});
    result = result | (input_112 & {4{sel[112]}});
    result = result | (input_113 & {4{sel[113]}});
    result = result | (input_114 & {4{sel[114]}});
    result = result | (input_115 & {4{sel[115]}});
    result = result | (input_116 & {4{sel[116]}});
    result = result | (input_117 & {4{sel[117]}});
    result = result | (input_118 & {4{sel[118]}});
    result = result | (input_119 & {4{sel[119]}});
    result = result | (input_120 & {4{sel[120]}});
    result = result | (input_121 & {4{sel[121]}});
    result = result | (input_122 & {4{sel[122]}});
    result = result | (input_123 & {4{sel[123]}});
    result = result | (input_124 & {4{sel[124]}});
    result = result | (input_125 & {4{sel[125]}});
    result = result | (input_126 & {4{sel[126]}});
    result = result | (input_127 & {4{sel[127]}});
    result = result | (input_128 & {4{sel[128]}});
    result = result | (input_129 & {4{sel[129]}});
    MUX1HOT_v_4_130_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_4_2;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [3:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    MUX1HOT_v_4_4_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_5_2;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [4:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    MUX1HOT_v_4_5_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_64_2;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [63:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    result = result | (input_51 & {4{sel[51]}});
    result = result | (input_52 & {4{sel[52]}});
    result = result | (input_53 & {4{sel[53]}});
    result = result | (input_54 & {4{sel[54]}});
    result = result | (input_55 & {4{sel[55]}});
    result = result | (input_56 & {4{sel[56]}});
    result = result | (input_57 & {4{sel[57]}});
    result = result | (input_58 & {4{sel[58]}});
    result = result | (input_59 & {4{sel[59]}});
    result = result | (input_60 & {4{sel[60]}});
    result = result | (input_61 & {4{sel[61]}});
    result = result | (input_62 & {4{sel[62]}});
    result = result | (input_63 & {4{sel[63]}});
    MUX1HOT_v_4_64_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_66_2;
    input [3:0] input_65;
    input [3:0] input_64;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [65:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    result = result | (input_51 & {4{sel[51]}});
    result = result | (input_52 & {4{sel[52]}});
    result = result | (input_53 & {4{sel[53]}});
    result = result | (input_54 & {4{sel[54]}});
    result = result | (input_55 & {4{sel[55]}});
    result = result | (input_56 & {4{sel[56]}});
    result = result | (input_57 & {4{sel[57]}});
    result = result | (input_58 & {4{sel[58]}});
    result = result | (input_59 & {4{sel[59]}});
    result = result | (input_60 & {4{sel[60]}});
    result = result | (input_61 & {4{sel[61]}});
    result = result | (input_62 & {4{sel[62]}});
    result = result | (input_63 & {4{sel[63]}});
    result = result | (input_64 & {4{sel[64]}});
    result = result | (input_65 & {4{sel[65]}});
    MUX1HOT_v_4_66_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_67_2;
    input [3:0] input_66;
    input [3:0] input_65;
    input [3:0] input_64;
    input [3:0] input_63;
    input [3:0] input_62;
    input [3:0] input_61;
    input [3:0] input_60;
    input [3:0] input_59;
    input [3:0] input_58;
    input [3:0] input_57;
    input [3:0] input_56;
    input [3:0] input_55;
    input [3:0] input_54;
    input [3:0] input_53;
    input [3:0] input_52;
    input [3:0] input_51;
    input [3:0] input_50;
    input [3:0] input_49;
    input [3:0] input_48;
    input [3:0] input_47;
    input [3:0] input_46;
    input [3:0] input_45;
    input [3:0] input_44;
    input [3:0] input_43;
    input [3:0] input_42;
    input [3:0] input_41;
    input [3:0] input_40;
    input [3:0] input_39;
    input [3:0] input_38;
    input [3:0] input_37;
    input [3:0] input_36;
    input [3:0] input_35;
    input [3:0] input_34;
    input [3:0] input_33;
    input [3:0] input_32;
    input [3:0] input_31;
    input [3:0] input_30;
    input [3:0] input_29;
    input [3:0] input_28;
    input [3:0] input_27;
    input [3:0] input_26;
    input [3:0] input_25;
    input [3:0] input_24;
    input [3:0] input_23;
    input [3:0] input_22;
    input [3:0] input_21;
    input [3:0] input_20;
    input [3:0] input_19;
    input [3:0] input_18;
    input [3:0] input_17;
    input [3:0] input_16;
    input [3:0] input_15;
    input [3:0] input_14;
    input [3:0] input_13;
    input [3:0] input_12;
    input [3:0] input_11;
    input [3:0] input_10;
    input [3:0] input_9;
    input [3:0] input_8;
    input [3:0] input_7;
    input [3:0] input_6;
    input [3:0] input_5;
    input [3:0] input_4;
    input [3:0] input_3;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [66:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | (input_1 & {4{sel[1]}});
    result = result | (input_2 & {4{sel[2]}});
    result = result | (input_3 & {4{sel[3]}});
    result = result | (input_4 & {4{sel[4]}});
    result = result | (input_5 & {4{sel[5]}});
    result = result | (input_6 & {4{sel[6]}});
    result = result | (input_7 & {4{sel[7]}});
    result = result | (input_8 & {4{sel[8]}});
    result = result | (input_9 & {4{sel[9]}});
    result = result | (input_10 & {4{sel[10]}});
    result = result | (input_11 & {4{sel[11]}});
    result = result | (input_12 & {4{sel[12]}});
    result = result | (input_13 & {4{sel[13]}});
    result = result | (input_14 & {4{sel[14]}});
    result = result | (input_15 & {4{sel[15]}});
    result = result | (input_16 & {4{sel[16]}});
    result = result | (input_17 & {4{sel[17]}});
    result = result | (input_18 & {4{sel[18]}});
    result = result | (input_19 & {4{sel[19]}});
    result = result | (input_20 & {4{sel[20]}});
    result = result | (input_21 & {4{sel[21]}});
    result = result | (input_22 & {4{sel[22]}});
    result = result | (input_23 & {4{sel[23]}});
    result = result | (input_24 & {4{sel[24]}});
    result = result | (input_25 & {4{sel[25]}});
    result = result | (input_26 & {4{sel[26]}});
    result = result | (input_27 & {4{sel[27]}});
    result = result | (input_28 & {4{sel[28]}});
    result = result | (input_29 & {4{sel[29]}});
    result = result | (input_30 & {4{sel[30]}});
    result = result | (input_31 & {4{sel[31]}});
    result = result | (input_32 & {4{sel[32]}});
    result = result | (input_33 & {4{sel[33]}});
    result = result | (input_34 & {4{sel[34]}});
    result = result | (input_35 & {4{sel[35]}});
    result = result | (input_36 & {4{sel[36]}});
    result = result | (input_37 & {4{sel[37]}});
    result = result | (input_38 & {4{sel[38]}});
    result = result | (input_39 & {4{sel[39]}});
    result = result | (input_40 & {4{sel[40]}});
    result = result | (input_41 & {4{sel[41]}});
    result = result | (input_42 & {4{sel[42]}});
    result = result | (input_43 & {4{sel[43]}});
    result = result | (input_44 & {4{sel[44]}});
    result = result | (input_45 & {4{sel[45]}});
    result = result | (input_46 & {4{sel[46]}});
    result = result | (input_47 & {4{sel[47]}});
    result = result | (input_48 & {4{sel[48]}});
    result = result | (input_49 & {4{sel[49]}});
    result = result | (input_50 & {4{sel[50]}});
    result = result | (input_51 & {4{sel[51]}});
    result = result | (input_52 & {4{sel[52]}});
    result = result | (input_53 & {4{sel[53]}});
    result = result | (input_54 & {4{sel[54]}});
    result = result | (input_55 & {4{sel[55]}});
    result = result | (input_56 & {4{sel[56]}});
    result = result | (input_57 & {4{sel[57]}});
    result = result | (input_58 & {4{sel[58]}});
    result = result | (input_59 & {4{sel[59]}});
    result = result | (input_60 & {4{sel[60]}});
    result = result | (input_61 & {4{sel[61]}});
    result = result | (input_62 & {4{sel[62]}});
    result = result | (input_63 & {4{sel[63]}});
    result = result | (input_64 & {4{sel[64]}});
    result = result | (input_65 & {4{sel[65]}});
    result = result | (input_66 & {4{sel[66]}});
    MUX1HOT_v_4_67_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_129_2;
    input [4:0] input_128;
    input [4:0] input_127;
    input [4:0] input_126;
    input [4:0] input_125;
    input [4:0] input_124;
    input [4:0] input_123;
    input [4:0] input_122;
    input [4:0] input_121;
    input [4:0] input_120;
    input [4:0] input_119;
    input [4:0] input_118;
    input [4:0] input_117;
    input [4:0] input_116;
    input [4:0] input_115;
    input [4:0] input_114;
    input [4:0] input_113;
    input [4:0] input_112;
    input [4:0] input_111;
    input [4:0] input_110;
    input [4:0] input_109;
    input [4:0] input_108;
    input [4:0] input_107;
    input [4:0] input_106;
    input [4:0] input_105;
    input [4:0] input_104;
    input [4:0] input_103;
    input [4:0] input_102;
    input [4:0] input_101;
    input [4:0] input_100;
    input [4:0] input_99;
    input [4:0] input_98;
    input [4:0] input_97;
    input [4:0] input_96;
    input [4:0] input_95;
    input [4:0] input_94;
    input [4:0] input_93;
    input [4:0] input_92;
    input [4:0] input_91;
    input [4:0] input_90;
    input [4:0] input_89;
    input [4:0] input_88;
    input [4:0] input_87;
    input [4:0] input_86;
    input [4:0] input_85;
    input [4:0] input_84;
    input [4:0] input_83;
    input [4:0] input_82;
    input [4:0] input_81;
    input [4:0] input_80;
    input [4:0] input_79;
    input [4:0] input_78;
    input [4:0] input_77;
    input [4:0] input_76;
    input [4:0] input_75;
    input [4:0] input_74;
    input [4:0] input_73;
    input [4:0] input_72;
    input [4:0] input_71;
    input [4:0] input_70;
    input [4:0] input_69;
    input [4:0] input_68;
    input [4:0] input_67;
    input [4:0] input_66;
    input [4:0] input_65;
    input [4:0] input_64;
    input [4:0] input_63;
    input [4:0] input_62;
    input [4:0] input_61;
    input [4:0] input_60;
    input [4:0] input_59;
    input [4:0] input_58;
    input [4:0] input_57;
    input [4:0] input_56;
    input [4:0] input_55;
    input [4:0] input_54;
    input [4:0] input_53;
    input [4:0] input_52;
    input [4:0] input_51;
    input [4:0] input_50;
    input [4:0] input_49;
    input [4:0] input_48;
    input [4:0] input_47;
    input [4:0] input_46;
    input [4:0] input_45;
    input [4:0] input_44;
    input [4:0] input_43;
    input [4:0] input_42;
    input [4:0] input_41;
    input [4:0] input_40;
    input [4:0] input_39;
    input [4:0] input_38;
    input [4:0] input_37;
    input [4:0] input_36;
    input [4:0] input_35;
    input [4:0] input_34;
    input [4:0] input_33;
    input [4:0] input_32;
    input [4:0] input_31;
    input [4:0] input_30;
    input [4:0] input_29;
    input [4:0] input_28;
    input [4:0] input_27;
    input [4:0] input_26;
    input [4:0] input_25;
    input [4:0] input_24;
    input [4:0] input_23;
    input [4:0] input_22;
    input [4:0] input_21;
    input [4:0] input_20;
    input [4:0] input_19;
    input [4:0] input_18;
    input [4:0] input_17;
    input [4:0] input_16;
    input [4:0] input_15;
    input [4:0] input_14;
    input [4:0] input_13;
    input [4:0] input_12;
    input [4:0] input_11;
    input [4:0] input_10;
    input [4:0] input_9;
    input [4:0] input_8;
    input [4:0] input_7;
    input [4:0] input_6;
    input [4:0] input_5;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [128:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    result = result | (input_5 & {5{sel[5]}});
    result = result | (input_6 & {5{sel[6]}});
    result = result | (input_7 & {5{sel[7]}});
    result = result | (input_8 & {5{sel[8]}});
    result = result | (input_9 & {5{sel[9]}});
    result = result | (input_10 & {5{sel[10]}});
    result = result | (input_11 & {5{sel[11]}});
    result = result | (input_12 & {5{sel[12]}});
    result = result | (input_13 & {5{sel[13]}});
    result = result | (input_14 & {5{sel[14]}});
    result = result | (input_15 & {5{sel[15]}});
    result = result | (input_16 & {5{sel[16]}});
    result = result | (input_17 & {5{sel[17]}});
    result = result | (input_18 & {5{sel[18]}});
    result = result | (input_19 & {5{sel[19]}});
    result = result | (input_20 & {5{sel[20]}});
    result = result | (input_21 & {5{sel[21]}});
    result = result | (input_22 & {5{sel[22]}});
    result = result | (input_23 & {5{sel[23]}});
    result = result | (input_24 & {5{sel[24]}});
    result = result | (input_25 & {5{sel[25]}});
    result = result | (input_26 & {5{sel[26]}});
    result = result | (input_27 & {5{sel[27]}});
    result = result | (input_28 & {5{sel[28]}});
    result = result | (input_29 & {5{sel[29]}});
    result = result | (input_30 & {5{sel[30]}});
    result = result | (input_31 & {5{sel[31]}});
    result = result | (input_32 & {5{sel[32]}});
    result = result | (input_33 & {5{sel[33]}});
    result = result | (input_34 & {5{sel[34]}});
    result = result | (input_35 & {5{sel[35]}});
    result = result | (input_36 & {5{sel[36]}});
    result = result | (input_37 & {5{sel[37]}});
    result = result | (input_38 & {5{sel[38]}});
    result = result | (input_39 & {5{sel[39]}});
    result = result | (input_40 & {5{sel[40]}});
    result = result | (input_41 & {5{sel[41]}});
    result = result | (input_42 & {5{sel[42]}});
    result = result | (input_43 & {5{sel[43]}});
    result = result | (input_44 & {5{sel[44]}});
    result = result | (input_45 & {5{sel[45]}});
    result = result | (input_46 & {5{sel[46]}});
    result = result | (input_47 & {5{sel[47]}});
    result = result | (input_48 & {5{sel[48]}});
    result = result | (input_49 & {5{sel[49]}});
    result = result | (input_50 & {5{sel[50]}});
    result = result | (input_51 & {5{sel[51]}});
    result = result | (input_52 & {5{sel[52]}});
    result = result | (input_53 & {5{sel[53]}});
    result = result | (input_54 & {5{sel[54]}});
    result = result | (input_55 & {5{sel[55]}});
    result = result | (input_56 & {5{sel[56]}});
    result = result | (input_57 & {5{sel[57]}});
    result = result | (input_58 & {5{sel[58]}});
    result = result | (input_59 & {5{sel[59]}});
    result = result | (input_60 & {5{sel[60]}});
    result = result | (input_61 & {5{sel[61]}});
    result = result | (input_62 & {5{sel[62]}});
    result = result | (input_63 & {5{sel[63]}});
    result = result | (input_64 & {5{sel[64]}});
    result = result | (input_65 & {5{sel[65]}});
    result = result | (input_66 & {5{sel[66]}});
    result = result | (input_67 & {5{sel[67]}});
    result = result | (input_68 & {5{sel[68]}});
    result = result | (input_69 & {5{sel[69]}});
    result = result | (input_70 & {5{sel[70]}});
    result = result | (input_71 & {5{sel[71]}});
    result = result | (input_72 & {5{sel[72]}});
    result = result | (input_73 & {5{sel[73]}});
    result = result | (input_74 & {5{sel[74]}});
    result = result | (input_75 & {5{sel[75]}});
    result = result | (input_76 & {5{sel[76]}});
    result = result | (input_77 & {5{sel[77]}});
    result = result | (input_78 & {5{sel[78]}});
    result = result | (input_79 & {5{sel[79]}});
    result = result | (input_80 & {5{sel[80]}});
    result = result | (input_81 & {5{sel[81]}});
    result = result | (input_82 & {5{sel[82]}});
    result = result | (input_83 & {5{sel[83]}});
    result = result | (input_84 & {5{sel[84]}});
    result = result | (input_85 & {5{sel[85]}});
    result = result | (input_86 & {5{sel[86]}});
    result = result | (input_87 & {5{sel[87]}});
    result = result | (input_88 & {5{sel[88]}});
    result = result | (input_89 & {5{sel[89]}});
    result = result | (input_90 & {5{sel[90]}});
    result = result | (input_91 & {5{sel[91]}});
    result = result | (input_92 & {5{sel[92]}});
    result = result | (input_93 & {5{sel[93]}});
    result = result | (input_94 & {5{sel[94]}});
    result = result | (input_95 & {5{sel[95]}});
    result = result | (input_96 & {5{sel[96]}});
    result = result | (input_97 & {5{sel[97]}});
    result = result | (input_98 & {5{sel[98]}});
    result = result | (input_99 & {5{sel[99]}});
    result = result | (input_100 & {5{sel[100]}});
    result = result | (input_101 & {5{sel[101]}});
    result = result | (input_102 & {5{sel[102]}});
    result = result | (input_103 & {5{sel[103]}});
    result = result | (input_104 & {5{sel[104]}});
    result = result | (input_105 & {5{sel[105]}});
    result = result | (input_106 & {5{sel[106]}});
    result = result | (input_107 & {5{sel[107]}});
    result = result | (input_108 & {5{sel[108]}});
    result = result | (input_109 & {5{sel[109]}});
    result = result | (input_110 & {5{sel[110]}});
    result = result | (input_111 & {5{sel[111]}});
    result = result | (input_112 & {5{sel[112]}});
    result = result | (input_113 & {5{sel[113]}});
    result = result | (input_114 & {5{sel[114]}});
    result = result | (input_115 & {5{sel[115]}});
    result = result | (input_116 & {5{sel[116]}});
    result = result | (input_117 & {5{sel[117]}});
    result = result | (input_118 & {5{sel[118]}});
    result = result | (input_119 & {5{sel[119]}});
    result = result | (input_120 & {5{sel[120]}});
    result = result | (input_121 & {5{sel[121]}});
    result = result | (input_122 & {5{sel[122]}});
    result = result | (input_123 & {5{sel[123]}});
    result = result | (input_124 & {5{sel[124]}});
    result = result | (input_125 & {5{sel[125]}});
    result = result | (input_126 & {5{sel[126]}});
    result = result | (input_127 & {5{sel[127]}});
    result = result | (input_128 & {5{sel[128]}});
    MUX1HOT_v_5_129_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_3_2;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [2:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    MUX1HOT_v_5_3_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_4_2;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [3:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    MUX1HOT_v_5_4_2 = result;
  end
  endfunction


  function automatic [4:0] MUX1HOT_v_5_5_2;
    input [4:0] input_4;
    input [4:0] input_3;
    input [4:0] input_2;
    input [4:0] input_1;
    input [4:0] input_0;
    input [4:0] sel;
    reg [4:0] result;
  begin
    result = input_0 & {5{sel[0]}};
    result = result | (input_1 & {5{sel[1]}});
    result = result | (input_2 & {5{sel[2]}});
    result = result | (input_3 & {5{sel[3]}});
    result = result | (input_4 & {5{sel[4]}});
    MUX1HOT_v_5_5_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_3_2;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [2:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    MUX1HOT_v_7_3_2 = result;
  end
  endfunction


  function automatic [6:0] MUX1HOT_v_7_5_2;
    input [6:0] input_4;
    input [6:0] input_3;
    input [6:0] input_2;
    input [6:0] input_1;
    input [6:0] input_0;
    input [4:0] sel;
    reg [6:0] result;
  begin
    result = input_0 & {7{sel[0]}};
    result = result | (input_1 & {7{sel[1]}});
    result = result | (input_2 & {7{sel[2]}});
    result = result | (input_3 & {7{sel[3]}});
    result = result | (input_4 & {7{sel[4]}});
    MUX1HOT_v_7_5_2 = result;
  end
  endfunction


  function automatic  MUX_s_1_2_2;
    input  input_0;
    input  input_1;
    input  sel;
    reg  result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [10:0] MUX_v_11_2_2;
    input [10:0] input_0;
    input [10:0] input_1;
    input  sel;
    reg [10:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_11_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input  sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input  sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input  sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input  sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input  sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input  sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input  sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [6:0] readslicef_8_7_1;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 1;
    readslicef_8_7_1 = tmp[6:0];
  end
  endfunction


  function automatic [4:0] signext_5_4;
    input [3:0] vector;
  begin
    signext_5_4= {{1{vector[3]}}, vector};
  end
  endfunction


  function automatic [6:0] signext_7_4;
    input [3:0] vector;
  begin
    signext_7_4= {{3{vector[3]}}, vector};
  end
  endfunction


  function automatic [5:0] conv_s2s_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2s_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [6:0] conv_s2s_6_7 ;
    input [5:0]  vector ;
  begin
    conv_s2s_6_7 = {vector[5], vector};
  end
  endfunction


  function automatic [5:0] conv_s2u_5_6 ;
    input [4:0]  vector ;
  begin
    conv_s2u_5_6 = {vector[4], vector};
  end
  endfunction


  function automatic [7:0] conv_s2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2u_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [11:0] conv_s2u_11_12 ;
    input [10:0]  vector ;
  begin
    conv_s2u_11_12 = {vector[10], vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_4_7 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_7 = {{3{1'b0}}, vector};
  end
  endfunction


  function automatic [6:0] conv_u2s_5_7 ;
    input [4:0]  vector ;
  begin
    conv_u2s_5_7 = {{2{1'b0}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    fir
// ------------------------------------------------------------------


module fir (
  clk, rst, input_m_rsc_dat, input_m_triosy_lz, input_e_rsc_dat, input_e_triosy_lz,
      taps_m_rsc_dat, taps_m_triosy_lz, taps_e_rsc_dat, taps_e_triosy_lz, return_m_rsc_dat,
      return_m_triosy_lz, return_e_rsc_dat, return_e_triosy_lz
);
  input clk;
  input rst;
  input [10:0] input_m_rsc_dat;
  output input_m_triosy_lz;
  input [4:0] input_e_rsc_dat;
  output input_e_triosy_lz;
  input [703:0] taps_m_rsc_dat;
  output taps_m_triosy_lz;
  input [319:0] taps_e_rsc_dat;
  output taps_e_triosy_lz;
  output [10:0] return_m_rsc_dat;
  output return_m_triosy_lz;
  output [4:0] return_e_rsc_dat;
  output return_e_triosy_lz;


  // Interconnect Declarations
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_1_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_1_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_2_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_2_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_3_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_3_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_4_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_4_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_5_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_5_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_6_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_6_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_7_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_7_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_8_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_8_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_9_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_9_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_10_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_10_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_11_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_11_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_12_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_12_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_13_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_13_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_14_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_14_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_15_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_15_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_16_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_16_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_17_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_17_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_18_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_18_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_19_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_19_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_20_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_20_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_21_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_21_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_22_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_22_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_23_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_23_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_24_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_24_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_25_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_25_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_26_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_26_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_27_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_27_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_28_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_28_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_29_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_29_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_30_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_30_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_31_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_31_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_32_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_32_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_33_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_33_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_34_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_34_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_35_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_35_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_36_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_36_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_37_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_37_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_38_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_38_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_39_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_39_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_40_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_40_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_41_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_41_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_42_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_42_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_43_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_43_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_44_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_44_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_45_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_45_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_46_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_46_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_47_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_47_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_48_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_48_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_49_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_49_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_50_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_50_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_51_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_51_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_52_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_52_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_53_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_53_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_54_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_54_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_55_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_55_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_56_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_56_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_57_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_57_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_58_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_58_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_59_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_59_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_60_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_60_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_61_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_61_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_62_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_62_rtn;
  wire [17:0] MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa;
  wire MAC_1_leading_sign_18_1_1_0_cmp_63_all_same;
  wire [4:0] MAC_1_leading_sign_18_1_1_0_cmp_63_rtn;


  // Interconnect Declarations for Component Instantiations 
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_1 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_2 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_3 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_4 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_5 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_6 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_7 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_8 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_9 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_10 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_11 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_12 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_13 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_14 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_15 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_16 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_17 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_18 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_19 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_20 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_21 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_22 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_23 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_24 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_25 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_26 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_27 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_28 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_29 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_30 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_31 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_32 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_33 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_34 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_35 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_36 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_37 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_38 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_39 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_40 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_41 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_42 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_43 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_44 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_45 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_46 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_47 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_48 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_49 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_50 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_51 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_52 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_53 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_54 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_55 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_56 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_57 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_58 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_59 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_60 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_61 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_62 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn)
    );
  leading_sign_18_1_1_0  MAC_1_leading_sign_18_1_1_0_cmp_63 (
      .mantissa(MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa),
      .all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn)
    );
  fir_core fir_core_inst (
      .clk(clk),
      .rst(rst),
      .input_m_rsc_dat(input_m_rsc_dat),
      .input_m_triosy_lz(input_m_triosy_lz),
      .input_e_rsc_dat(input_e_rsc_dat),
      .input_e_triosy_lz(input_e_triosy_lz),
      .taps_m_rsc_dat(taps_m_rsc_dat),
      .taps_m_triosy_lz(taps_m_triosy_lz),
      .taps_e_rsc_dat(taps_e_rsc_dat),
      .taps_e_triosy_lz(taps_e_triosy_lz),
      .return_m_rsc_dat(return_m_rsc_dat),
      .return_m_triosy_lz(return_m_triosy_lz),
      .return_e_rsc_dat(return_e_rsc_dat),
      .return_e_triosy_lz(return_e_triosy_lz),
      .MAC_1_leading_sign_18_1_1_0_cmp_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_all_same(MAC_1_leading_sign_18_1_1_0_cmp_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_rtn(MAC_1_leading_sign_18_1_1_0_cmp_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_1_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_all_same(MAC_1_leading_sign_18_1_1_0_cmp_1_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_1_rtn(MAC_1_leading_sign_18_1_1_0_cmp_1_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_2_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_all_same(MAC_1_leading_sign_18_1_1_0_cmp_2_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_2_rtn(MAC_1_leading_sign_18_1_1_0_cmp_2_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_3_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_all_same(MAC_1_leading_sign_18_1_1_0_cmp_3_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_3_rtn(MAC_1_leading_sign_18_1_1_0_cmp_3_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_4_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_all_same(MAC_1_leading_sign_18_1_1_0_cmp_4_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_4_rtn(MAC_1_leading_sign_18_1_1_0_cmp_4_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_5_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_all_same(MAC_1_leading_sign_18_1_1_0_cmp_5_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_5_rtn(MAC_1_leading_sign_18_1_1_0_cmp_5_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_6_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_all_same(MAC_1_leading_sign_18_1_1_0_cmp_6_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_6_rtn(MAC_1_leading_sign_18_1_1_0_cmp_6_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_7_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_all_same(MAC_1_leading_sign_18_1_1_0_cmp_7_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_7_rtn(MAC_1_leading_sign_18_1_1_0_cmp_7_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_8_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_all_same(MAC_1_leading_sign_18_1_1_0_cmp_8_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_8_rtn(MAC_1_leading_sign_18_1_1_0_cmp_8_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_9_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_all_same(MAC_1_leading_sign_18_1_1_0_cmp_9_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_9_rtn(MAC_1_leading_sign_18_1_1_0_cmp_9_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_10_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_all_same(MAC_1_leading_sign_18_1_1_0_cmp_10_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_10_rtn(MAC_1_leading_sign_18_1_1_0_cmp_10_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_11_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_all_same(MAC_1_leading_sign_18_1_1_0_cmp_11_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_11_rtn(MAC_1_leading_sign_18_1_1_0_cmp_11_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_12_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_all_same(MAC_1_leading_sign_18_1_1_0_cmp_12_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_12_rtn(MAC_1_leading_sign_18_1_1_0_cmp_12_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_13_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_all_same(MAC_1_leading_sign_18_1_1_0_cmp_13_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_13_rtn(MAC_1_leading_sign_18_1_1_0_cmp_13_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_14_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_all_same(MAC_1_leading_sign_18_1_1_0_cmp_14_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_14_rtn(MAC_1_leading_sign_18_1_1_0_cmp_14_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_15_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_all_same(MAC_1_leading_sign_18_1_1_0_cmp_15_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_15_rtn(MAC_1_leading_sign_18_1_1_0_cmp_15_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_16_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_all_same(MAC_1_leading_sign_18_1_1_0_cmp_16_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_16_rtn(MAC_1_leading_sign_18_1_1_0_cmp_16_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_17_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_all_same(MAC_1_leading_sign_18_1_1_0_cmp_17_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_17_rtn(MAC_1_leading_sign_18_1_1_0_cmp_17_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_18_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_all_same(MAC_1_leading_sign_18_1_1_0_cmp_18_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_18_rtn(MAC_1_leading_sign_18_1_1_0_cmp_18_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_19_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_all_same(MAC_1_leading_sign_18_1_1_0_cmp_19_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_19_rtn(MAC_1_leading_sign_18_1_1_0_cmp_19_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_20_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_all_same(MAC_1_leading_sign_18_1_1_0_cmp_20_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_20_rtn(MAC_1_leading_sign_18_1_1_0_cmp_20_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_21_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_all_same(MAC_1_leading_sign_18_1_1_0_cmp_21_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_21_rtn(MAC_1_leading_sign_18_1_1_0_cmp_21_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_22_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_all_same(MAC_1_leading_sign_18_1_1_0_cmp_22_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_22_rtn(MAC_1_leading_sign_18_1_1_0_cmp_22_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_23_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_all_same(MAC_1_leading_sign_18_1_1_0_cmp_23_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_23_rtn(MAC_1_leading_sign_18_1_1_0_cmp_23_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_24_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_all_same(MAC_1_leading_sign_18_1_1_0_cmp_24_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_24_rtn(MAC_1_leading_sign_18_1_1_0_cmp_24_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_25_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_all_same(MAC_1_leading_sign_18_1_1_0_cmp_25_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_25_rtn(MAC_1_leading_sign_18_1_1_0_cmp_25_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_26_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_all_same(MAC_1_leading_sign_18_1_1_0_cmp_26_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_26_rtn(MAC_1_leading_sign_18_1_1_0_cmp_26_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_27_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_all_same(MAC_1_leading_sign_18_1_1_0_cmp_27_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_27_rtn(MAC_1_leading_sign_18_1_1_0_cmp_27_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_28_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_all_same(MAC_1_leading_sign_18_1_1_0_cmp_28_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_28_rtn(MAC_1_leading_sign_18_1_1_0_cmp_28_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_29_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_all_same(MAC_1_leading_sign_18_1_1_0_cmp_29_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_29_rtn(MAC_1_leading_sign_18_1_1_0_cmp_29_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_30_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_all_same(MAC_1_leading_sign_18_1_1_0_cmp_30_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_30_rtn(MAC_1_leading_sign_18_1_1_0_cmp_30_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_31_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_all_same(MAC_1_leading_sign_18_1_1_0_cmp_31_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_31_rtn(MAC_1_leading_sign_18_1_1_0_cmp_31_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_32_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_all_same(MAC_1_leading_sign_18_1_1_0_cmp_32_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_32_rtn(MAC_1_leading_sign_18_1_1_0_cmp_32_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_33_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_all_same(MAC_1_leading_sign_18_1_1_0_cmp_33_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_33_rtn(MAC_1_leading_sign_18_1_1_0_cmp_33_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_34_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_all_same(MAC_1_leading_sign_18_1_1_0_cmp_34_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_34_rtn(MAC_1_leading_sign_18_1_1_0_cmp_34_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_35_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_all_same(MAC_1_leading_sign_18_1_1_0_cmp_35_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_35_rtn(MAC_1_leading_sign_18_1_1_0_cmp_35_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_36_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_all_same(MAC_1_leading_sign_18_1_1_0_cmp_36_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_36_rtn(MAC_1_leading_sign_18_1_1_0_cmp_36_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_37_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_all_same(MAC_1_leading_sign_18_1_1_0_cmp_37_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_37_rtn(MAC_1_leading_sign_18_1_1_0_cmp_37_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_38_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_all_same(MAC_1_leading_sign_18_1_1_0_cmp_38_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_38_rtn(MAC_1_leading_sign_18_1_1_0_cmp_38_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_39_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_all_same(MAC_1_leading_sign_18_1_1_0_cmp_39_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_39_rtn(MAC_1_leading_sign_18_1_1_0_cmp_39_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_40_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_all_same(MAC_1_leading_sign_18_1_1_0_cmp_40_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_40_rtn(MAC_1_leading_sign_18_1_1_0_cmp_40_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_41_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_all_same(MAC_1_leading_sign_18_1_1_0_cmp_41_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_41_rtn(MAC_1_leading_sign_18_1_1_0_cmp_41_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_42_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_all_same(MAC_1_leading_sign_18_1_1_0_cmp_42_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_42_rtn(MAC_1_leading_sign_18_1_1_0_cmp_42_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_43_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_all_same(MAC_1_leading_sign_18_1_1_0_cmp_43_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_43_rtn(MAC_1_leading_sign_18_1_1_0_cmp_43_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_44_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_all_same(MAC_1_leading_sign_18_1_1_0_cmp_44_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_44_rtn(MAC_1_leading_sign_18_1_1_0_cmp_44_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_45_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_all_same(MAC_1_leading_sign_18_1_1_0_cmp_45_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_45_rtn(MAC_1_leading_sign_18_1_1_0_cmp_45_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_46_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_all_same(MAC_1_leading_sign_18_1_1_0_cmp_46_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_46_rtn(MAC_1_leading_sign_18_1_1_0_cmp_46_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_47_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_all_same(MAC_1_leading_sign_18_1_1_0_cmp_47_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_47_rtn(MAC_1_leading_sign_18_1_1_0_cmp_47_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_48_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_all_same(MAC_1_leading_sign_18_1_1_0_cmp_48_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_48_rtn(MAC_1_leading_sign_18_1_1_0_cmp_48_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_49_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_all_same(MAC_1_leading_sign_18_1_1_0_cmp_49_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_49_rtn(MAC_1_leading_sign_18_1_1_0_cmp_49_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_50_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_all_same(MAC_1_leading_sign_18_1_1_0_cmp_50_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_50_rtn(MAC_1_leading_sign_18_1_1_0_cmp_50_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_51_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_all_same(MAC_1_leading_sign_18_1_1_0_cmp_51_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_51_rtn(MAC_1_leading_sign_18_1_1_0_cmp_51_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_52_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_all_same(MAC_1_leading_sign_18_1_1_0_cmp_52_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_52_rtn(MAC_1_leading_sign_18_1_1_0_cmp_52_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_53_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_all_same(MAC_1_leading_sign_18_1_1_0_cmp_53_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_53_rtn(MAC_1_leading_sign_18_1_1_0_cmp_53_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_54_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_all_same(MAC_1_leading_sign_18_1_1_0_cmp_54_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_54_rtn(MAC_1_leading_sign_18_1_1_0_cmp_54_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_55_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_all_same(MAC_1_leading_sign_18_1_1_0_cmp_55_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_55_rtn(MAC_1_leading_sign_18_1_1_0_cmp_55_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_56_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_all_same(MAC_1_leading_sign_18_1_1_0_cmp_56_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_56_rtn(MAC_1_leading_sign_18_1_1_0_cmp_56_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_57_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_all_same(MAC_1_leading_sign_18_1_1_0_cmp_57_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_57_rtn(MAC_1_leading_sign_18_1_1_0_cmp_57_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_58_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_all_same(MAC_1_leading_sign_18_1_1_0_cmp_58_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_58_rtn(MAC_1_leading_sign_18_1_1_0_cmp_58_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_59_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_all_same(MAC_1_leading_sign_18_1_1_0_cmp_59_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_59_rtn(MAC_1_leading_sign_18_1_1_0_cmp_59_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_60_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_all_same(MAC_1_leading_sign_18_1_1_0_cmp_60_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_60_rtn(MAC_1_leading_sign_18_1_1_0_cmp_60_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_61_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_all_same(MAC_1_leading_sign_18_1_1_0_cmp_61_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_61_rtn(MAC_1_leading_sign_18_1_1_0_cmp_61_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_62_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_all_same(MAC_1_leading_sign_18_1_1_0_cmp_62_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_62_rtn(MAC_1_leading_sign_18_1_1_0_cmp_62_rtn),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa(MAC_1_leading_sign_18_1_1_0_cmp_63_mantissa),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_all_same(MAC_1_leading_sign_18_1_1_0_cmp_63_all_same),
      .MAC_1_leading_sign_18_1_1_0_cmp_63_rtn(MAC_1_leading_sign_18_1_1_0_cmp_63_rtn)
    );
endmodule



